PK   �rZrr���=  ��    cirkitFile.json�}k�%���_��b��a�L�7�3�k���`��$\�sT;����j�^A�}ɼU����&��	Uc��[UI�<�|D�t�X���?����/�ㇻ�����no�����ߪۛ�w�����<�￿y�S��x����h��kb�C�uT�Q�n}(�LQ5]]�u�q��?���y�����������C���UY����EUֺ0�����*o����������vu��v.�:�3	���,�wg�Q�µ�*lW�E�{_4M45%������w�����b������82�e���"����Q��l��-C.�:�l\u�L���Q��ͩ8jI���������!�4F�ـ����G��]B�y�4˵��h~�O���gS��9h�X�������ɟ��d	�;�L^�J�M͙h,i�.F%��Ǩ�ǁ�p�����EP�<�L\��>|&.�E>�A]r�39p�%�7�A]�W39p�E�3�H,%�T�m�%W/�o�% g�K�^.!��z������mߐ3�� mZ`C<{�L����SB�u6��@���G�����,��"� 8�|oZ�m:B�u6�G���������vj��dC����f����o;�*m�_��4|�Ɇ�,���Y �"����m'"���N6Dd���l�Ȃo;���v�!"��dC����N6Dd���l�Ȃo;���v�!"�B.�vZ��dCD|�Ɇ�,���Y�m'"���N6�:8��dCD|�Ɇ�,���Y�m'"���N6Dd���NǷ�l�Ȃo;���v�!"��dC�Cɷ�l�Ȃo;���v� ����1 \ڻ���a٩aeGX�A���������Q�F!�Y�`p���[�+�Y�`p�[���X�A��]�_��sX�A��]�4��+����#,�ٍ���Lk�mcMzj���~����C�b����-�������-�	. GS`����c���� �
8�#p���G`~�[<�%b�.��Et��w�x��ų�h�Y ۼ�9�������y�px�#��kv{���k4Y����;��#� ���� d���_�E���>_U�7���hBe
k�.j�7�	��#eu�\=#p�h�iLQ������؃/ϛ��,�d����Af/`[��q��������]U����=��s�17��+�uFX�!~�b�JMe��ì��X~旮����(F���~���� ���X~�X~�ˏ���D���۾X~���� �����Q����]-*��"�Q��Ɔ�xуcW,�tI,?p���G`~�z/X~��V,?�K���3�V,?�KW���G=X~�.����z���/]c�}�}��p�c�Q�����`���,?�KI���.X~��5���?���/%� �`��_J��8���#0���+?�?���/�%�`��_J��8���#0��
,?p���G`~)�X~�v�v��Â��?���/%�`��_Jy�8���[�z*]]�&Bhj��*EE�b�*��P��c �6-�y��`��������j/���L����J��ժ����.�*���wZ�P�5S��M��A&w���ή���4ZhST�Xˁc-,?�K	����ZX~�Rǁ������/%��ka��_J��:�	:�	8�r�Xˁc-,?�K)���ZX~旒;������/����`��_J���_	����#0��
,?p���G`~)�)X~��ˏ6���*�4�����Os��>M����4������;�OsK�>M
���4�����4�{Ն�vL��}to}��;q��>S�fr�[��}��?�ޟ��|Mr����8���x�j�a��8�&֫5�՚�j�y5��-W�x-w��$^�Kf�yo�����\�6I3���<�6�V��+S����~�5h��
74}a���}�hꪵa�=��C�S���u����f�uὋ��Ml|Tѵ��j�2������u;�}�bh�_V5M�LD��>4��e��oϪ��vE�+��(�H>�]Q�!�]�DKV����gU_{��\6��f����9� �AEs�L�Z��@[�J�E�T�I�;o����Q��z��y:�NƫyN�����j��E�eƫYNօ'�Ֆ�����r����3�qΫ�4<��zM�3�Ϋ�ܺ�W��Y��c����!{�,^ҫ�*��Iez �Ae}+o�;��̚6gMq�W���)����1�5�q^�6UdNq�W���S��k�|ߖ��n0ѯ��E�B4{�ZS�mm/9�Y��]���1MV���V�Qo����
[[Tm��Q��'���cΨ������mϪ����4�*Cu�UN7EPM�]�zҥo�������mϪ������m��j��E�����M(��t4�v�����VV�:�S����T_o{�]�wT���6U_�U�n|�U���R۳�_��rY��iZ-nh<M�Ơ���)�T�ʅ�'�暪�:z]��E��A���Z�C]_��Y��55��8J���û�Ǜ�?�V�����WJ���z B�V��Wj��c'��_��w|F �q������#��W��Ȣ9��@@*E�F ��q=�f{�*U�S��U(F%��bD�����k"���D0�M�����T��a�LN0�M��¼ ��F!��� g�tQ♾�� �@@9�[&#г��`���r� �m�]�[�(F��6�� �Ѷە{"�h���dRnW&#��p�2��T�וk"qVg�av;����y�r���#U�׿Yur9���	�	f�QH/��̂̄���x��	f�	f�QHj<r,av\��8
I�G�A�`���q�߃8��p��($5�q��q��($5�q��q��($5^  ��0;n`v��>j�[I�-��츁�qR���̎�G!���0N0;n`v����8�츅�qRJd���f�QH)�6�nM�(��f�QH)�2�̎[�G!�̾0N0;nav���K��~`v���8
)%�q��q��(�� �	����ބ�q��(���	f�̎��R?'�/av�����8��x	��kH���Os�Q�LpT�J"\�a���
��W�Ӝ�K��,T�\�\��@�Ns�c�:ͨ����+(�i�u8*P�\I�k�D�:�����W�}�N3�c$ ��D���4W;ƾN3�/���/�9W�\�\r��p��>s���p��	Ls�c�u��#�9W0*2.�	�H&�aK2l��f�%��K(쒉�H"�9�E�V"L$�鬹���D_lѰH��`$����%�|?1�����yd��j�Bd+��L 6�ւ��L(��"�`l�~%[�pl�-D�� "[�(�dؒ�t7FF��H��2a��t�G���y����[Zb��f����Dؒ�t�JF�B;bB[b2q���t�a�����Dئ;p2����Dؒ[u�)[��1���(?A&.�2;dl���t�RF��ɰ%�鎨�le�2�$�6�u����n�[�a������엉�%��le�2�$�6ݡ���L\&dئ��2�:�(t\Q&.32q����Dؒ�t7_F�2q�[�a�r��V&.aK2lS����e"lI�m�� #[��L�-ɰM�+dd+���%�)��l�L\&dئ\"2����Dؒ۔EF�2q�[�a�r���V&.aK2lS��
�$�J&�Y�����e"lI�m�$#[��L�-ɰU����"e+q�dئN2����D��[����ݠs�V&.[`��Eދ��˦�6�caKKl!B��˜L\&dئg2����Dؒ۔�MF�2q�[�a�r���V&.aK2lS�<�
e�J�!�9�����e"lI�m�e(#[��L�-ɰM9ed+���%�)���le�2�$�6���m)�_&dئ\�2����Dؒ۔�TF�2q�[�c�>���᾿:�m?P_���-,y_Te��I���v�;�;QVr��DY�&�e%��N����;QVre�DY�n�e%�N���;QVr>��:��b�w��{a0����ֽ0^���^�?Z�N)ˁ����[��{��!���Fc`f��*I��?���,���T� �9~�p�����mq��P�����P�CESW����6^M
���@T[3غ��E��&
&���Pu�m��ݢ,���vh�0���ƿ�j��I�+�!\YV��撅��EE����"�5�(�]Q�!�]�ԥ��z�K�&��ŒM��5�el�����M�TE��S�d����N��/ПǶT�*�ʩs��/���@����E��6�آaP��(c�3���2�KCSv�g�ؗ�I����J��ժ���e(�*���wZ�P���ğ��9�g�lN�Y(��~ʦ뚅�9�g�l:�Y(~k4f�T[�!e3��ӺMc�C[&Fo��<�ec�`양Ƀq[V����m
�����.D���Ck꺭m�l���9Cf�l�BY(���7Q�YO���-�6��Ѯ����Y�uʦ\�P6咅�)��4�*Cu��N7EPM(�kZO���S�r�BٔKʦ\�P6�R7����6h�k}�PM�hp���U�Ji��8�A�G9(�r	�k����S�8٦�ສЍ��*4}Sf�%e;о錵E�hL��k�7�	��#e�s4pi��B����P4�l��Tա���.Z�>� ���Ժ�:��e�l�Qʩ��<�������O�aO>GWuQ}ȨB�>��EU��E_�������r����w���
�h!�@@G�
a:Zg#��#�c#��"#�c,#��5#�c?#�:Ƒ���8���3�($u�1�`��`�����<��~̀g e�����e@@9�[&#P�������A1�����P���m�P#Р���2m�]��@@9�[&#P�������H��ƙm����r9�,w�ו�	f�3��\N0��u�r��o�ׅ��f�QH�x��	f�	f�QH�x
�X�츆�q�:���p��q��($u<�����f�QH�x��	f�5̎����+�̎k�G!��9\L8��f�QH)�=�n%����f�QH)�8�̎�G!���0N0;n`v��2)�8�츅�qR�����f�QH)S,�nM�(��f�QH)�'�̎[�G!��0N0;nav��2¶~`v���8
)eȃq��q��(����	����ބ�q��(��9�	f�̎��R�&'�/av��2�8��x	��kH���̲H�Q��x �$D���,�(W	�$�Uf٣Ш@�Jp%��0��F�U�+�p�q��\g�|!��J"\�$"�Y"_�$���裈�u��"	�$�Uf|Ѩ@�Jp%��0�ދF�U�+�pU�Y�^4*P�\I�k:,�D\"lI�m:�,#[��K(쒉�H&�"��K�-ɰMg�ed+}��%��̼�le"0�$�6�����L&dئ;2����Dؒ�tCF�2ј[�a����V&"aK2l����De"lI�m��#�� ���%�鮒�le�2�$�6ݹ���Ў�Ж�L\�e�2-���%����le�2�$�6�哑�L\&dئ;�2����Dؒ�t�RF�2q�[�a����V&.aK2l�]W���e"lI�m��+s0I&.aK2l��c���e"lI�m�C-#[��L�-ɰMw�ed+tZQ踢L\fd�2#���%��n��le�2�$�6����L\&dئ\	2����Dؒ۔�AF�2q�[�a�rW��V&.aK2lS�Z��L�-ɰM�Ddd+���%�)'��le�2�$�6�v���L\&dئ52��I&t�L&.�2q����Dؒ۔3HF�2q�[�a�r��V&.aK2lS'���e"lI�m�E%#[��L�-ɰM9�Dd�d�2�$�6����L\&dئg2����Dؒ۔�MF�2q�[�a�r���V&.aK2lS�<�
e�J�!�9�����e"lI�m�e(#[��L�-ɰM9ed+���%�)���le�2�$�6���m)���%�)ק�le�2�$�6�,���L\&�ض?����}��WeA�oK�UY��h�C�;��]��N��ܴ;QV���DY��e%��N��\�;QV�[�DY�G�e%��N����{����]���^���}Zu/F��>`���k�	���ⵏq��`�k��}Xr/F��>߸��kI����O�����9�pC��ۡ�����Zۓm2����ET[3غ��E��&
&���Pu�m��ݢ,���vh�0���ƿ�j��I�+�!\YV��撅��EE����"�5�(�]Q�!�]�ԥ��z�K�&��ŒM��5�el�����M�TE��S�d�`�d��T�*�ʩs��/���@���(�EY(3S
�E�R��Tunp�m�jUXM�2�A^S�;�U�Ͷt�P6����)�,�M�f�`��9�g�lN�Y(�3~�感��9��iHy1ڻ{��`�w;�ʃ����:߷e(�L��R�]����붶�u�f?e�lvS�f/��zY��T��آj����Iy�5[g�l�%eS.Y(��kK����n�j��"�&�5�']�֩�Y)e{\�l��M��M5�F��E�Z_�&�ES:\;�u��R���=�rP��Qʦ\��ھ���T4N���"��*t��
Mߔr�Bَ�o:cmф*Z=���Ma��;�HY��`�l�Q�v��j��^�t�2�q(�����P��.eS.Y(�r��6��_��û���]�כ�F���x��8�WG�9�������7�0v�<�����6<O��j��8�&�7�y����+�Ό�XK��W�<w���5�]o�zep�.�s^�y[����*�d��<����ۢaq�^?�p�<*�4�*�Ge����
.��u*a
��69���VeiS�oɢ2́ɡBL*8�W,p�sˑgڹ�b�m(r�	V^��������G�N���:$�r9��u��ȓ�*t�Ca�`���ꢯCh�SuP��i���_�P2M����KGM���Z澞9�N��åC�P�`�+�ݛ���v¾}���G�h��J�^�_�+qd����|;_�L+Q�6�% ��F�碒����a΅Fp.��A��K��~2���G<O_4T2L2H&�2�犂����p�Ͷ��ۖV���g�/:��,kel�5�eM��-��M깯���Ϯ�si��V2����׾�z�˕�t�գ+�pv����^|�}����G�忖�|a�w�}�ݲ��{`�������6C�� pǄ�0w�6�|?\���0u���jv�r�OAy�<*Q*߽�z�x�K���n��7�t,����_�l�������������E���=>�)>>�a>>�>>��>>#�	�����������K���l�
'}i1E�%^��W9��g�>��Y�Л/�E��G/2x��|F背�^�g\`�k��nİ@r|�����̩��J,Pa�}}����g^�x�c������\5�m�_/�y~I�;�{��_lO]wlx���`JO$<���]�<W��$�W_����!�0R"�5�A̽��N�C�Z��s�r19�v���+�`��W'�@$ ���Q'�n�/gX3�+�U'��Ț��DN��9q�q@ý�X�\��X���	�M�מ��/��
�!�\p�~�� �=�D��n�]��z��V��������F�ˈ��_�Ͽ�q�ܥ���^�A�B0��� )�;b���[j����Cb:�%�KR`+�����Y�����oƿ_Й�u�,r<�/���u	H����tq���t �2/_j%�B�Q�-��ޫ�2F�'|���D~���]7�ZF�AI~�r�E��+_���b{����������ۛ�����������(������]w��'�~��u�ǘ�ј�;C���ǿ�,\����&�b�%D�8×B�ܜ���HY>)�B���d�`C�����Ľ �����ְΕш�$�b?��I�L,��/!��h.,�'�ݦ3�:"CGH.-3�S�	`�in�5W� ����1Ƌ���qukr�#�t�/����qً���,.���L|�j&6���U��U糸43Y�!.;f�,���ɂ�.�M�,�ꢣ�ɂ�.;F�fa=�`?/�>���3�lͫξ7�5���Z<�K`b�'��e��h�.�.#�Rx /,/#�? x ��_>�J��<�+�{��`m�*]u�� ��`O�*] �� �S��|�R3�y ��S>�JW��q'���=�cD {�ǈ<� {j ���y �)#� �S>F���|��`O�)�-���Z�=�cD {�ǈ< ���y �)#�@����S>F���|��`O�����1R�y �=u {�ǈ< ���y �)#� �S>F���|���g��`O�����1"�=�cD {��P�`O�����1"�=�c�?�Ώ�#��!k&����:X~�����R�]>�̂��sF���'3���sF���n����E�,?����E/,�,?,?�%��|Հ}�t
��1cϔ�.S�X;�q2?f��Ks���ee~)1����.㙣CB�6`��f8϶|�R#Rx��x�造�n�d,CDh��L�/3��1F�=`��,AFKѡ��<'����o�]����cq� ��AKs�\C�K�$3��k	��Ӝ0W[�#[!����\	�����g�~��̿��%Lh��Fظr���>k��n�>Ϣ��Ӵ\�0aZ ̕ z�I�#/0CB3LWV�2��.���С��F.��c+0�tU-CtlfHh��Z��%0CZ`8���=i�nӜ�D��Є��3�H����a�8��!: 3$4�t�-C�f�!���`�v�!��˖h��0CB3LE�2DG1`��f�.��e??��b:�1�(̐���b��Q�!����h��0CB3L���2D�)`��f�.��e��S�	�0]�G����aJ ��E�)`��f���e��S�	�0%`@����aJ��!:N3$4Ô�-C�%�-t�b�q�E�)`��f���e��S�	�0%KA���N��1a�	��/h���0CZ`8�#�y0�q�L1[tP3'��#E5n�Ds��	�a��1�C�8`��f��"�e��q�	�0%tB���aJF��!:�3$4ÔH-Cx�x�t���1�C�8`��f���e��q�	�0%_C�Ԁ�aJ��!:l3$4Ô�,��fHh�)aZ��8̐�S�A��q
�!m1������ꫲ ӷ�%�ua4�ӝU�ο9���,a����D�;����?KT���,�����İ;����?Kĺ��,��^�a+ W���������p�p�}�� \=��/��śT����{���s���Ϳ�8����=*��3s<��>�h9xn��8x�/B���s<����͒�||h?3���/O� 4��P�����E=�P4u��0؞lsѱɩ�}��Y���f�uὋ�M@Tѵ��j�2������vh�0���ƿ�j���+�!\YV������ޯ��teu%���+*=����뚺�u]_zV��/],�D�ZS[F����'o�SŞL�9��y;d�����f�N���?�?mm�*U�S1��IY:o����Q��Rcժqɀ[��Vmi��Զj�2�f���Ȃ�Olj�+����m�]�
�)ڍ2��k�}��
�Yꊕy7.��Ȃ��2���bũʂ��Ggտ�Fgտ�Eg՟�j��d��]�h�P/O/��<�e^1Syxڼb����y�P��-��K��7���LUm���2�&��ϩ]�>Z���u[ۋ.BV�StV�.VV�q��7QrYO���-�6:�q6�=)�_\N��Ϫ��Y�/��2���PA]7D}�MT
�֓.}�ԥ�gտ����ڟU�B��z�u����/Bʢ)�����v�U����Կ��9�/�?���;��NE+b��/��B7����My��Y�/��7���hBǯ��~m��0���u����\�W)n>�Њ��7�\hŷɂ��-��y�Tա���.��>�~����P�mWV�}�U���?��|�w�����۟nrV	n�~s�&�4)��6M��!HZ��.	(�<9Q��3&Dsꍙ Ǆ��Ό==
t�1�#�1JWFt�1����l���c��1}�����>�n����Y#8��]����+�D�grB�
9��9q�r���9�����r<���bŜ)v�b�ܴX1Ǩ/V̱��j�a��ߔ1�'�m���п���?����Q�ծ��Y^�qذb��Fsذ"���pذ����r�p�e�6n�M��k?gΦ�Y]3������6���%��8lX;Gj�M�a~�dz�fƎ�ls�*����X֜ݹ=���iRi��)؜��ҝ��ѭ��~͢eFp,vӴ�svk.3 �s[]�6�sw�9�[36zmgnH�d5�]:g��qe���U=��=����z'_K��贓Q�n}�bPWTMW}Bc������,0:�zW�r?-�٣��P�Vgr�S�9.#�-ܖ�J.C�WM�C�e��fm1�������)�����ָ5�iYXS���s~Ĕ���1�)?V��
�#T.Z���N2fS���`�3GF�O�3���ë�0y���f4��Y�����sOv�k4�3Q��^��{��E3�Q���J��%&�
�v�m�[����[�{�*-�R�eX�2ܽ�:g��֕s����.�S�קû��ߥ�5�s���_����t0yBϏh�H??��G����?�Ϗ���{~����G���~�珪�G��Qx~f��E4�4��-���Ѽi��4���^�F���M���/<���~�6=�7�����_ڧ���/�������y��K���}�������K��y����\̋\�\.�E.f.�"3�����s�����\̋\�\.�E.f.�"3��yi�Yh����\f��>���>�\�<��xxy-�����߽;�L w�����݇�d.�B�����>�`�h�������cWK+����X7Лp���Cux�Oɘ�?M��~J��?������}��t׏�T~x��I�F�O�w�i&��H?���7��}L?�:uV�t���]l�M���?�����Fܛ�CjP|�����wͻ���������n�>Eⱓ��?u����D��	�������I�������(�o�*�hw������4���Z7�t����9Ux�ڢV���l�o��֦a�I���?~�������S}���N��<<�E����fT���}�?��7��o�*��ml�>��N����tؕ����b�)�?}� �>B������(�jTk5¤�y��I�\��V'?��O��p�Ĩ�'F�Y󟟘�b��<}� ����kO�}~0���d��%��`.���MOF�ҥq蜾�u���Oߎc�ۛ���|������ۛ�oo��7��j�P4��U���hL5����u݌������??����Ǻ�P9�*�m��Z�0�]An�,U�Uc����zCSahL��).��5�R�ŵ��hJk=|������N_�(I�b�U$lu4㽫��Y�C��2ݱ�~��}��c�ɷ/v�sK~��ݻ��+��7�P�}��:]4��EW�ޥ�P�+�D�������O������eG�}[��T���3�h��D孳K(�}��?e3�������N���N�~0��m���������>�K�3��>��ߤY�w���������ۏ�c�ӂ��%�O�~x|�u�=�><?���n�v��ݻ~A���=C?+X]Ry�)E����~����A��T}��Ú�3��7mQ��b�5�Vu�t�ʦՃSK
fO��]QW��:⢂��)Z��X�7��̸6Tm�&���(��TT���F��E�S��=����_>�O������O�~{��W��_��}������'_��_}�?��_==|������8����?���=<,��P��/�<����������������}Ufd�󭺽9Z�?�����L2�i��ϻ�??}��>M�7�Ƽ1Q3���?�'�w��E���?;'�>���[�j�'2�G�/H}��ӿ��g\�[p;.��q�������o��t����mm��Q��n��[�������S����?����vo|b������^z���DK\�u{|����.�� /�7�q"{��V�}c*Fe)ڕpK1�|c�sw�2C�{C������f���B_����v��T&���Te�8c�1���X0*����b�R�WV�|U�8����6xzC�26N���Q������ֻ��)�nmY�0�	������ն~d��ߡ���!*{�R������*R�h��*���&'�]���Q�]T�u�N�����;ﭏ���5#�B�.�A'��19)�5N�p�TrK.&Kʕ�L4UT�8��O֔ї���������:[��d�&�"HF|��ƞ��D�r�jTi�OP�QU�N��j��Ok�j|G�#��W��c���pc���̖�>?p�M�)ٹ�+J7�Ո��c@�WpC��Q��JR*��3+�zc#Te�sS�1�c嗦�?ה�k��r��F|s����4�G���)�s��sq���������p��_��w�l�o����귟'�0:I(��h��w=����/B���R�uS�B�Ъ���i��n^��٤�1*PUҘ�0�ӟ��9{��[���=��^	�UU
�Uֽ�=ju���o+�Y��kص���K@͂>j��r��˺Ι�o��X�����w������?��\}���t�s�w�-Ҩ,�까])s�m��R.�RJ��'�o�.�DI�?ME��.��(�`K*ʡkbP���ic��B�(��;�	��:���AEq���OeS�ONHyl��=S������1�Qm�w1�Jލ�m۩�����9W�3�+r�M�1@����7eY�3g��YN���3_��(�O�lA1�s&F0��Oљ�o�7���1C�&Ƭ��b ��iL]FI�ٲ���Ǵ�9+{B��2����lA�짣��O|a�����}ώL�
�w���/�l%�WA���xS4��?^5�Bm�����4"kЖGa����(�ZU��';��*'>��_���B6WN�U�����*i��ٲ*�W<�mt\�7*�X�� 1���L�B��ijh�NǮ��������,uN��i�?���
L�)�^V]\���/kZ�ka�1/��e&ڣ���ėN/=|��Ʈ}zx�R��z�Q'�ޤ��7U4�I?�uO�'���M��/����;uq4�Q�U)����~J�S����o>����z�ۿ��?���ã����7�=<�������qO1�������]��b7�ﻋXy�9F����?C�E���{�pw��u�����ӷ�~{�N��i�:=���~H�}�M��Ӣըm����'�M��<��>;�ϲ��R-+˫�}�����V��~������l�N�P��8�4h��P�4��䧅VQ'gŨz\4��R�T����t}d]�r��<e31J3Pe38e�he3Pe�W)ۧU�Y��%�se���F�x�EZ-(�v�3���E������g۶�*��)��MC���R��-��Ĳ-(۴؊�%˖Qly5�G�w㕋�;+�����6` �tR�u��:�����mS��S+:y6�e�&�g�,V�Er�l�b�ʦ�� �Me�ZV"4���|]˧�W��d�2�:բ�bi�d����mn�pj�>KG���Y(�K�d���J��6�X��nR~9]�/+۴�Z)v�E��T���{]��4y�k���u'�r'�Uw�;�Oo�꾜�r�UwZlE'ib��_j��d��*���K�;wbs��h�3YaR��Bn���<v���v/c>�w�lçŬ_.���if1e5�hwU���y���S���n|T]Au�9^���/�2��^�~9$��U���se\.6�2j�Zg���
DU��o,R�*�M����B+��+�x|��tyr{�@K�f����Q��Y5U�����Q�L�[�!S�e��א�F_�.�٪�Փ;�4V%��*���J,�3Wz����R1�~J^�o�L2~�O3;�;|���?��;�J��XK���-o���qn�LE����ek�*��ҟ���htيv<��
䦋��]�r�T�Yn>�=�W]Yn�T��W˜���������E���;��5�5�~<L{�U~٭��[^����U�V�Ny^1����o?@-��S`�X^��ݭ�˻���rˊF�_WNd���@V��+'�\�*�@w�
M����дܲ[G:\W.w��R�e+t͇P�S_�R�����"�>�'z"Wy|j:�,������4-F+��Y0���,X^U8Y^�i��+�0j[�#�e�l5����i9;��5/�X�J	X>uY�vIJ�ƌ�;N��ݩ2�U��	>K���h�ݚn�g[Y�9�S�]���<?�?�%��7,�߫�&o^6YK�>\g�d4����g�5�l�7y��[YbS�u��r9?�2����!CQ5���摀�-��j���R�[�,O{S�,���fo�*��z�j��x��Z�J�?*4��P-{�y���	��(����=��˄��=p}��S}[>J6Yn�+U-�~�5�����vQf����_��t�c�%S�u�_�Y��\��V�(��B�G�[ly���Bpf��5�X����%�7��`iE1���.S}ϋ��+"S�7��_^�:ϱ�Yj�bI�{�ES���r�[�7�<�^/��O�������K���/E�ؑ�RʙT�^`/6tYY&������7�2Ke�JU��Z�"��f~,Ƣ��|Y�"��jM��$�+F�7$���|^1u�����������:}��	4i$v\"�k)]u\b��e�;s�2K�Eu9��]LѢ*RW[�
��n���n�W�@��3f�5�ҝ��:$�K^���I�/�M�m^�jY���`�,��x�H���ϡ���"ϯ������맹�r�T?���=�*U-�v�z�SJ��E�3��lb�Y��4�L~���q����Y1���+T y�f<���p5C6���^���{�K��a�mC�#�8𷇧�bkK��b˛��;ߙ�py$X[�h����J@�#���y&f�+�5)f���+��)�2��,� �rw���n�l��e_�=�����i��m��#S���@؝Q*%�x�.[����+�t	4��Y^П���,T�+\m��ڗ���jo�]Đ��jOk��jO�/ϐ��+��>�r��ݟ�?�O��]����ۤ<���o�����X���������~�������ۧ�?��w�?Vs���PK   �}rZ�$&VAS }d /   images/6227b039-7cc5-4ac4-8a39-c32f35a7f912.png�PT_�/��� � �����A�9�d #9g%H�,9��0"9Ð$#�a�0C��3|߹瞺�^��[��U�]�k�{u��ի�ou/������S�caa)�Kkbaaoaa�cs��lq���N��XX���V���&@�t��w�r�t�|�b�����i�`��������Uڞ(�c,�W�^�;K��i<�B�Ր|b'%B�Q{]I�s�iJ�嫃\�oa���ͿVA^>@�����'O��U�Ka�t�z�0�5a�-�Zw�!Ȱ�^�~%��e%e��������9rֺ�m���6?`�/G</��6��>���%���~���#�y��7���%�_��%�L�U�<�Km�.P��&8&r+�ͼ�_��~d�N���a�c��v������ #vv���U��3�y����>�X��p�>V�6- Cr�O�ˁFo�/���n�*��v�v2Z�ny���3����hՐ����G�w>F�4w�bL$_%l���d��5��E���%�Ln��P�8����ܒO�]�&�m2�&�����'r�c[�����`������x���t��GX}i<�J�!��Z�?�>w�gÝ"翙zv�~�\_��^�3w��,![s@����-Fa	�_}1-�^��1j�ﻝ����}����-/,����jֹ�s��㲎��x\_���^P�5%+F�e��{C�������R�]=�=���N[:��8��mF�UY �	����P�9��R�&��f�.���Se➂\C��xn��>���٫H3h"7�}��p����6G����?
��f8���\&��ɿ�����U⫬ed�=�u��t(y ���a���L��n�v׭�^a䨑�6��� 4ت! ��W�ڝF��+g#��O�l��&��8�yk!u�W�]<�QF�r���@d:I���"h�n2mֵo ಑��~Fߑ�E�9~��b1^��Y��D�	gng@��[��$��/.������a��\�nW�u�w�>�b�?aۍ��-��1Iw�vs�A�,;�P�s��L�Y���o	xF$\KbwZBB��^&��6m٬)5��>�p��՜�T���N3�G�=��0�A��{����;g"��>��c������X�]�e
Z=ϋM?��?&�T�W	��3��!J���&�M����4�2��!j�k{+�B5N��},z�J~��/���e�V�t�X=�Y:� �\b�~-��2�������l���Q����̷Q�狨�����3��}���=G"���b2C$�)�k�� PH�X��4.�*.:�j�)����P�u_�Lißԡ�PԆ����cϑQ����V���n[�0�gt�r��&
��W��%����B���J������򙎶�\V��{��s��K���t�οs��2c��c�*����%��'b`����'�b�$��O�]�AeS>�i�l��=f���Ɖf��(l�̌m��;�_���D�q�I�߻�q��
�)�w��N[@v.�i�6;��J��k-�TnLd��V�<bҀ��#/�\�L�|d`V{��e���]����3~Ÿ�_O�0�j�uJ���܈j�gP��Bt.�n/�h���ƌF�����Y;���J�x��դ^����*�{�Q5�*ݚ��*�q�Q�v�J(G�D���ذKL;#f�Ni�N��s�? Y���2A��h�&��,�4��ֈ�ky�{�XqM�0��C���F-n�0��Q�#y�Dn3���x���N$��6X��1l��A��@��%GI�p��b����p�Ձ/��Q�)�
��͔k��쬇�O�삂ȋ�����4��
=�+���%�I�m����%wL	A�r�L�~c��h ����ѯ(UH�ců�h���=���v�TV7pE��Z�w��n?����&h���L��"�ƛ�l�������5�	gWa;�&��	gJ5N���ݶ�� ��5uʱ�}��lᙬ�٢5��Ǎs����8���\]$�ۣf�I.��'�����ƺ�*'������K�3����Dmf����51H[�f�6R��T�z����T��kP�R����U Ѕ�+U��K������uCGp��y�-����QG;�5�#��WO1n�b�Ą�mE��޶r��ά ̂���d�ap����Ӓ��j��)�}k n�Ep��%���K�J��Ք�;[�_�#uI`+��6]�(|Z<�\g�y�˧뒹a��;��mJ>N�Xν�S�kHlQ �$���``��l���Lb�D��L��L��(@�~�j~��*1,������arS�Y%����4i�*1w�q����7(v�$3Nd&\yr	�����r�����1[)�u0^?�Z�ġ�&=)� �ܴo�hy�th����J�����D#��ck�U�vq� �IvF��G��8> N�c���O�CWc�(T����㫑��-������o]y��:�f��Y��O��<w?d�}�	�	���sa�C������+!�Vf���R�[y��qF�g�� �+@ZC�+�;o`��2Ua[��2r��Z�:�Z�<���9 	p|�-�����8�_�/C��:LZ���T-v 
f����f���IY^�P�,���#`Mø����%^Ed�Ty6�@�{e&(	Q$��V��z42?b�D�N(��ƍ�V�I̔�[�pҌg�m�V�=K�F۬&�^_�T���9}�?Q r�?�y'��>�qW;��-`ǲ�=>��e\�������=(�'{�+��h�ꀝ�r�=*B��ȧ���{y �ENЛN%�$����+�&����@~�q�F�-$�xhd�S-�L����L
����+/�2u�?p���H�Uo�\�|E� �Qm��ȑ��fZ�l�eЁ��,Z��w\�웭�\k(�8���5(T�jd��u��Im%e�����2����=rsI۫�U�������9İ�$Kl#B�+�wn"�Fvx���TC�PU������	$|b���|rЊ���c�e� P��ܢ�>�x\�ì�^�+ Ϙ"��b���V�/�Kl��7\�p)R�����Onkŉ�G\��3):�j���7��J��\��/-�^Ƈߎ��u���N@���]D����l��r��X\�T,�Xj�QE���M*f�>/������_!��_�U����Zm��͊�WԹ�/��b���F/�s�ds)�fL��|���\>=#���Q!�<�=���>���h`bM×g�f�jf���,&��~��c�=+���Ą>�6.�h�c>�&���$8#���X~���+p���z�Py�g�1�\���|j�'Ծg��� ?�Nx�'��	.���1N�Ax���d��a��6�)�u�d�?^�x\�V҉ӄ5�{�,ik�=r�����չ��m�}Dq t�*�W4�Al����κ��Dں��k�2qľU%��6φ-��yѓL����ý�Ck�P�R�HC=c�TP���̣-lT�
�Òת�5oe��N�X7NJVI�o��F� X�n�%�@��R���s4p�S��H��1�)���> -H��W���2��j��u�{#�&����;�����v���5)%�s;�|�*����=�v�d�ts_���G�ux��Ү��qLw,��U��Yt��%�VX����"����������Va���6��adߵwN?#���\.��Z�
H��4�T޺��=I�=�yu5aڣYxu.0�u��p7vre0����B�!�2@kuc[��F������fނ�����D+?�o"�b��PjX��jG�hw���z���i������Zl�L��l�ᰢ/A�M����F��!|}\�7�s�{���.5�6U�iE��߄L�����-�g��3���j�X=$V�Gy�[��Q>�!�ӟ7x��}h��A�u���9�2���b�l������?�����wUGFņ����Tb%Z�u����C�s�(|�s/z0o�5b�|+h�d�s4��0U&ֿ�L���:��Ǆ;�b���we.��W�M�S8~�g�j3��x���;�����Xdz7���f~M��*�ōF�f��'`o��^�H��	�F�py`�\�o�<���IG�Lc���(46^~���n>�.��E�[!1�A'�ji�ɢ1��V��NNJ���C!�� VpMvI~D����H���=�ӨCx)�ɠSTe����4T���t���]ߚ�z�3L(,ml���fZUr,�HA=;_t�68o�?q�l��I0`�9)�Lk�8[������ "t�wr��~qcK���p<�P�������O>)��"�Ў6Ӟ�9H�*tS𚯵�ڔ�Ԉ�Vn��n[�B������a|���`n��.y�|rU3�����̩��������t�w?���h�ܮ>�����#f�yJ���&ʤ�������a�M�1�
����x1,�`ӒAY�^u��ͥU�Ԧ�:P�.�d�b˃�l���tи�m7c;�AB]a1�;�a	��
6	Q�6�C�E Z:_Ʌ COF��b�c��gk�r�Ǐ��L	dU�O�E]��!-j(^��W!+����7rΌ����?���Z��a���icMޣ������S�\E�M$�M �bO|�nVa��� �Y_����l"����D�D��dD7�቗�@�Sǚv p���������P����6i���}� "E�騳�l~�k��W���d/�$�Y|z&�f��������R�-v��-7t��Z��|mQ�_��u�>%�4�u�C>=#d�;���CZ��WW�'KJ�<�J�gQn\=-�c�
 E)�H�5ym0�p���`�&Dm�zX_�|��y�1iL��]�B��U6��v:h�lk2�#��L3�v5gXrv����?s��k���"R,���f���2�2����#�p�5�LZX��=��H��e[лR5;b��Ig#����#݇��3Q ��;k~�s��� c�Ap�%>���j���nƕ,�l�J.?�[�t.�I����֦4�~T`��	�Ewo3'-���� r�;����� �Ze@���S@a{< ��� ȳ1�#r(U���[X4k�"J�D��$>qDq����9�e�K��ՠ�M���$E������.����G>e�@S���Ji�sl@怮�k�z��h2Ť4G~��5���� �7���z@���͑1�~��0M�	8NԷC;R��	��1�Q�" �:m~u{GWF���:��枯�0�j���8�\S�����(W��l��R�!X��f���[����t���i�th�<��}C:�?X�%G�z�<^S��	�J!kH8i斳�s�n?E�&V^�XN��zi�i�Vؤ�M��}���u���!�>GVJW� á1����uH��Ew� �he�:2h��(K�OJ=�a?�]f�_�k�Kw�7d'�lS陹A���٤�����@c�����$f�9HM^�1Q��1	�1��!�\�5���6�ن��F��O1J���|��S��3���#u��/	���C�=;ށ�~�j�D-��%G�M�JW���-����W�*�=P��#���N���I��2)	�Z�x�]���#\�/��dbZ �����o�/n�e�S�Gn�I��g���n�At����Ԕ�w�BX�_��
"���W���U�!��]�,á�n���u����o����z��/��蚸�m|ϐ234��k|���4�$%��Y�ȮFӂ������(��Kff�tB\c��R!5��q�-��~;�'����鐰*��>��~,����E�H���y��,��r�$KTT��������ؒ����bB�͗�����;���Cأ��mm���kwc��N"�F�i�g�KM��Pf��)W�f�򠖲!"��yw�K�&p)�_N��Ѥ������?W��`){b��Ƃ4������LW��(Q�������`N�ŝxm���v�!��{�Qt�l6v�!= �Gޖˌb�n�tſsu�d���ꮠ���Q�/a�+��={�s<�T���	ș�6�  Jh�L+-�.qOG��������w3��֠��iP�'������ �y�0T��ڱe���l)~����g��w��cc��ȶZ𕖲�����-Ty��b������&*
�Ќ:�r%�f����>Q���V�7V#�2��6]eA9M�U7`�QVOxG^ -�􎹧8S�"|�DI�hȕ��ï��������I�vZ(�f+��¤$�3�9�>k��:+@���<�*�P	�doZWf*q���l
	=9��W�+�_q�6��#@�@����(w��h�����ۅ�x��͛hU����z��/�+>�kce��;*�P��\�i��/'�K)>����d*+�Y2�([ʃ�_<��)K�֬dq�����	��I�}'��=%!X8QSS�27�^�U��=�X��5�{�-i�w
�^�xA#��@��g�c���r̾M37iͶ�M�>'�*J����(�k�<YE@�"SzZ듵rP�RcИ��b�r�{�Wb��D}��Wg�J���F!�VF�x�� �;����V�v��wfػ�|�sW�@��B�`ƛ}|�K�r4�RȨ)��UI���(���������GC��9)**�A�%��w�#2��_`���w����9z���/�{;҃S^ptFG�@�@�2�Z�����Y0��dU׳Q���+i֜Q>�Co��K�?�({�jҗ����U8�D��9���FzϴG��3ɢ�Z�N!�
W��.54�<�I�`�E����{[�
&�&��ܻ�/'�ݬk�q�%�Q�!	�7��*KJdI�m��6z�@�y�I�f��)R8 ����įzܐBsCY:����n,'}�5?�h�_w�H4�/�9=�]��CG�M�nt@��)/��r~����͸M��ĴK뮁V^ ����Z&�(�.�mh�,}A����-�+¯�e$"6sL���%��s�«W�2(�t+��n�v
�����W�uI?�f�pb9���O(�C3�(�m�e
��jl���M�e|���ߛ��X.���a_�\Ӓ@��"d���G��oI�f��Si�ּ�SPFY�+m&"��ak]�����T
�]�p�ׂ>��g��
�y����a�ejat�S�'��Ή浿�� է��w����=�ȏ+9��㢊�o��-�<����hl\_qStz�-�Fԯ]�,� �F1�qn�4���%ci�f�������F.�<���JT��NŮ��k��,�iE�����[���}u��Ϫ}6��1k�s����s���e����i�ÚN��CXp��HN㐽��d�U�a��И�1�$}�XD,2�
���p�4�
�@<�����m� (����T��P�VB��� �N��n��V-{�x�I���r����I1��t:p=]!&V��2!p�='���g�i���Y����v����1��iv�"���|N�u��V������[@�u;p�����VP<{��d�@�� ���*qQ�(9tݎ��PϺԽ�VVu(+��ǜقtB��4�c������=�zY����Uu%�qR-��N�Y���yX�P��"�{G6�C*�ס�Ֆ�~97�c�a
Z
]Ӟ��jZ�P���*�����I)6��7��`��T~�T�2����K�$b\Q����Nm� ,� ���;٬�,��a`}1B�<��5ˎ	-��E��	���~1_=ty2F�lj̢W�&��W@�-�Ӥ���xmt+6���y�(��2[z�œ�C�ZLaU"�/�'�je�D"9���b��m6�V��h�����m�o�RI���� ���k���?Sm���ъ��� T@A���� ��%�e���>ɛI?B+�JVI_~���aƕ��z�F֢��������?��B݀UY�Jhs�[�ۗno���7�ҭ�dP�!������9oL0mƨVtWe�럪����&?&�&�?Y�&J	;C�
�?��J{)�`B�#h��LÈ�6�S~L.}A�7nU��W�klf�)�]oJ�
�#]��Ų ({�?�w��1y�b7�	�7:b��Q2XHN��YԿ@Ar ��"^ �k�@H��\@g���?=cX�>���k!�5�8�@(i�' x~��2O_h�������Ԁ91/)g��{�<�l� $�K4�Pǧ3�(�s`�`߽AnH���D"���T�0��\}�\� �KH忛8�˽R�.��0�i�8��=��l��T�[��!M%^r��KSE:�e�������!
 X�����x� �&$����{r"�a�h[���2Q*���7�����1{��Z
[�:4(8��a�.�ihR��P�һ�d��p�?�կP[8=A�j�X<g��*�NV��{F��<�L��?�7sz�=˲�F۔���x;'^����D�C������f�vV�� �'���j��s �P?��	} gP'����'
�T"U_Õ�����t���)���r>��k���o���]�=6�S%��4�d����Ĺ!�"�����HrŹ����ۊ�Ŋ���z��&�d��w0���gI�j�( �1g����[�h��4�8N�͆^���޸�A�Fτa��~��[	�Y)�Ex닺+'��l��v^��D����#��V�ɳʠ���/1��f�]���m��R��B��(� 5�Z6C����aM�[9a������G�176�qW�t��7I����JaD@� �I�e�z[��LO_:w("��J���bJ����V��2�^�|�C��ߔ��Ň{�՚ƙ+�����EMʝ1�,J����ʌ����,:���mi?}V�D������&�pЬo$%�;���B��k�8պ�gG-�C��7ܯ�B/��H��C��(�i�gQ�9��/�ϠZ�Ǵ|�Q����������Ґ���%��Y�l
��b�]Y�{0y,ٙz��h�*toǈ%�`�JX���TqE���)�Ҕ���߲�I��.�{�>�9�7~?���V����i���^�l;�M��(��ة�ft��.S$X��M�b�̝1�^K�db�J#���J��/�wƸ3�$�O9.��͐���f�d?,�3c��N��ZuӜ�/�V��+��ή����t53�oq�]�~Ӷ2��@Y�N+�W�]��6�5���UE�J�U�Jq�����[�>��t�Y�Ѓy��0�ei�H�^4�ӊ���J&.������_\���m��^��@TD)q�nM^���N�R�W���A��Ӆ��ˡ\��yz��h�%"��� ��ǵ�Ac���v�3��y��Nx�-�T��_fс�w����<�,�Y�R$L�|�Q��[�2��A��#�;���G����|ٳ9�0��gԯuK�%M+���8	�X�_�hLzWm8$N��V$�Y/��|��w4�Np)�~Q����%(�^���܅>�{Vr���%������iL�0��]?�3�L���W����p���!u�{�w�-��I5����&��YT����F��
G�3�8�|�,`�r���G�r�����V��m<2�{*��X�p���g�P�a�f��w�5�4k�~tH�,@��@R􇿹m	8�2]n\|^Fl��޻�	@fv�LO����Q���W�y�X���Lg>���~F�Ô�WJ��и(x�� Xi񿜒��=8�|�@�]Q>N6O�
S�����GM���a�'����"dL�\��?�֝--����|�]���ԅ����m��Y�2m���=��P�r�OLǾ4�vQȊ�y#R��~����@M��@��g�C�1d�9���9kq�6������L��O���yS�5A���6>���@��G�5㽩�������;g^���c�c�u�8�av�8�|&ze㑀�ې����[�Bo����r�q���}V)��j*pN��Lx}���|�+�����n:C�ϓ��I�tF�Bh��ְ΍�le�V(�?h���3^�coʍ7�ؗ:V��eI+/����@[�����'N�8X{�C�SB�������������}9�`��?,>zs8���'FAus�hvE���ÎC���sn�-&��R:��G3�I�%��h玿g��nV<�ڮ�E�+��&۴ZMva��~p�n����ĺֿjR�E�1ʹ0v/X�ӷq��ح�L�5�[�l64L~�3fچ�}K~�����%�|	��?b�aHe�R����}t �B��[H^{����Ӏ�!zH���t{��i�A��s��yo�[�7�s�����x�Z�^���0� Z�&��R�-���䂌�W���ͷ��mg?�h�#���=�C�{�Ƒ������:�/�*��N�#7�I]��I���9�*�X�a��AT~5�*� �㿵���<�%�q����Q$\[>�Ê�
M����e�ݮ/�~"�'
'9h����Xd�Px�L�-}�p�����zj�� �\|�o�V�7d��>c3y���9��S
-�Fx�*��t��>)hyQlt�s}`S״��O9ΐZd|ѵajX(��(�C~*?���{*kZv���9��~�~k��U�����/���`�b�ې0��G����/�K_@d�CT��GS�B���%ƫ�/��^>G!�K�>��1��w���E��P�C�2:5w�V�{?N�������.d~E����ljY\9z`Ԥl�U�of�`n������u� ���^��fЩyl���k^�\��,H����ջ~��[M����	��+��[��:BP���[5����wuI�vc]҄�E��M�C�g=���?��R��3H���L��2u?�3'u����A�ep�	*n3�CLwI�v3t�/��h�Q�vM
q�J��yT�,�)8E^,�p��/��)��7����������ՙIBw�eb��'̼U�RC�ӆe�˼4�р ��l�
)�h�\��)���t
�41a������!�E'�(°ҟ(-u���U��%���i^�j.�����Hz�̍呂:YgD��?��̚��7�+Ϻ�9=��)���V�u`hx�G��Wb����{=�'K[3��_�� �������=z78ީ����Π���V$�ŻE?�Q"�U��?�N��k��WC�l�$eR��o�	���|�@BYW.^��I+��tK�nB��a�G�%#�=3�g��8��CF�*v�����u�P�ČE�9̄b']U�䄝��#3���u�gDJ�s[�ĺ
Z�|����[*E����f��+�������Y22��ƥ�yX�$�P�%m�i��N{���ғ!�*�����Ͱ�����݊�����P-h����Fidg�ݿ�>���F�Ϥ�6X�FNES��Ig��bW0�v ���𶢁�������Q��{6 �,.$Z5�͏5��k��NS}��1w�s���M֨g'B��!�vs��ݏ�
��.�����q���@.�N�j`W���t|5�*��yQ�����~��@?i>��^�lTd�}��6��Ҹ%��j��ϯ�~|淽���0�11��M),���r�����bT�()	���Rm�y+��Ӭ�������Sg6 \4�&�Fs��}�,I��a��՝�vs�;/��Ϝ�d(�>���_�뢁����m���')��@���fN���#�[
�G���b�M��NH&la`W_G�@%����<<_ro��"ˇ��L2xF�\O� ��﭂��z�S�[�_�]�K��c�����$�]��O�(֌���8�]=�����e؅���K�ȷօɯk4t�͜}x�d��:���u��������6v(S����V��M������ù��'�mp����f+9Έ� ;�ee�!D��ffUּ��22��F������������zk���(j-���ʞ�/��Zͅ&������J��M�CУ��jmw�KK�y��X�����h��������f�Y�{{�::��EEt�����-�EǻE|v3͜!.$w���@r��t��I-Dffflg+M��<������������*�h�U{���k}��4_gCEM�y�D�����u����i�@G�5�5-�8���j<��C��|�[�Xd|=:�c�1���Ղ2�r�]N��7�n��>�_����4С�����#G���ֶ��~턾<�JK������r?�4~{H�� �p�EHkkk����k5�k�������+r���
�XO[=v~�DQ$��1�����!���Km�v]!D��9Ӈ痀�f tT��[/��[��wf�;.�s5�����jYYv�����U����l���:dS#fM�E
T-��RI@`+�q�Ĭ�:��a�J謀P �B���� ܂�jUv�S�ɣ�e��C��>�%.�WZV��C�αk�`H����u4�X�U�4"�:���u�W-jj�fKM4�1�t��ΐ�(�9R%f���(����c�g|��9����}wϲr���]�:<-��zEU����])VK�Ik ��<�`�[3;��׍�lqcJ׷.���^�yW���ol�,H�� ���3YDG`Fր��UTj�d����An��}�9ꢸn�V�"H^E�~��k̕��@�$���QK����Ş��CO����Mv>j��R����Gww��{��tta��D@Is̀�b�@U����Q�HH�
���fJ��/�=��4�H���J��y���ʋ@���o�Vu{�]�gYi9�Ʌno�/Ɗ�&�+�-��#�he�s�NtO���,���#��Qﳞ�p\,	�A4^��u�g�G��Bz{>Q.�(�"��ӕP��i��#|5c��8|�0e��M Z���w��T�!\:�x�г�]��a�tvƈB�5n�R)�Y���1T]��r�������Пy���6���:	�	k����������-��E��iu�t?{�W�F8�2PE�����,�iz��!��4�h�����:�֋����D�WF��t���������!r�| #Y>��Zl�wPD�ɢ��F�i�s/�	��܎C�*k讃i�Q�JӲd����\`����V`��kk��#AW�EEV{X&2��ߎ�����J�Q��(�\	"�(0�|�"1_v�ٜ���0�������j0��H:Q���G�D.2��I��t�:+�HO�;g�"K��sRóp�I��@�[j���Z���NO�@�7�
�L�	�ȍ�H�����.��\M�5�"� ����>HJ�����l��Q�RJ�����)��=�Ԓ��Â���.�$[ޫ�����s��,������9�b�}�a��|�9����O�� �GK�`�(��W�|�{��:���.�#�c��v�Ň7�֫�\�/���ږi-�H�[���5|�K��N���ƪ�^����9��Y���mU&kl�=�뜙���~{�r{��itpn�w����	C`tW�3SS	�RN�pP�Ѷ���TuoJ�LjZ��ZҨm�Mp����Я���Y��eÇ��=ۙ4���R325�y���QJXD��$����Wm��q:76,.\:V]�	�����PɮRw�bN�B�R�n%7	����&!��:<��=��c�a�������>c�&��2�I��������=�=Gb��(@�̰�<+
��]����<�J}�K��5�S����~��7�O߱�IVU�����2�|���e�\��;bOظ�n
��
�-q)��:s ���^�7�q�p������E&6���.�*��xJ�	vvs�a= i���s�Z�S��j�f}�?�S���K�L�;����et�g.IV�C���6�
��2~��r�_"�lՇ(��6���u%3���Q��l����P��q�_n�]Z�B�w�+ C����Q�qE"Lˆ� �V|��'�����D�����w~���D��a w�y6x�L�NM�a��J�jn)w�[������cN�M��51s��S�h�9 ��z0��o"-�_I,J�!��@����c�����]X�i������� sy�LJ��w�f���3�z���O�]��b��r}�R71,���%O/m�+���Œ�*��p��!�5��������^�ĹgE��'�B���I[[cC���_otZ���N�����3{�|0c���o�ϴ�̟�#Eŉ�y\��Hr�����000�A5bˤ���F&X	���i�m~�|[3o�\8[ov�r��5O̫QZ�$�-	^��[1��a��	T^�P8f��>	����2�M�۲�^���r��Y_��XD�.ya��2q��L���]����U=�^�P��5Bd��X�a��.f��,ƞf�B{�׮h�D������Q)���_3����g]�tI��ZVt�et�����%zd������R�Ԟ;��o.�m� �S%T@f3���̎~���_�V���#�hx�z���ޖ���~�;[��{�ڻz�
�yk$���������GJ~P�)z���n%��W� ��qe@_����%�
���3���p`/���o���5���q��Y"�R�t��l�j��w�p/�քSP��b���	W����wf���q<�x���m�IU}�ƑoU|������:H��ҏ���2���9���ŭX�ۨ��.��D��N��N�Ғ��G�Yy��8]B7su_0r�C�3�'p�z6
�����/�O��Z
�n<B� 0"? 7���z��1�\���%��1Ά�\�lO~a?�W+��r����]��6�����^K��v/`,�&)��~������~|1C��̼:T�Fl�Qr�Û����j����V=0{T����Ȃ���� ��Q�E�����A˻�N��t2E�g���?O�����I��oz8VZl#���]��:Yl������C���>M9ʂ�::#��5��m8]�l!7V�w�m=�t�aJo*-'z|�6�����!��	AhQ��H`���cO��QJKK��ٍ����������7�Z"&��ߍ�yh|U�Yr��.���r�ӯ]��#���x�|��޽{4��M~�%(--}��]u�G��;a��d�>N�~�� kbbR��xG��K�Wlʖ�?5P�]�IK����Ib_�FRFߛ���;�v-y������r���j��f�W�_�����K\��fff��г��ٚ�޵�G/��M%�������}o����i�Z�IVzz������Z
^��dլR����_5Y ���`F��S�@3i���;s�E��ܣ�
�}��f3���~P�kkOm�++)u��|�����We�^*�Y`\�U���}�OP4�]����W�/��%�I����;��1�c8]\]�W��ؠ!Du�ll�Sp��}8����$��̃XL��!���F��U2��o��D2�Y�5���RL�үܕ�r����=n�3����{�}o��叏4��q�[m����a)<Vnͦ��amK�n´���ʪ:B�:P�З�m��oZ�l���~p]�L�/��-��8�%qx]��}��ߡ�e*TI	�����Z�	%3��X����3�$&,���b7sW%M����������e��1"�� __���ѯZ�]\���:�׼�adaY����|u}?�}�Bă}mm�b��~�m��!�8�0��}��� 凕�1y�ʲ鯩��Ŀ�p���>�|΋(W듖��������\\\�!.���N w��&o�F|Ğt�fx��qv]_�G����"`|00w8Z�ͪ��{w�7��|�S�۹��*y�c�݆��A��w��g&���8�v3��G����N�ڲ��✖�g�F|�5�%3jrЪ�������R����ᖴt��XA��^����$F�p�H_�~�����h``�n���+Q���Z)����o-AG�<�u�*��,õ�<V�pcD_Tv�X����ᝓjQ�GXy[�EEuJ�}���Hz����{���������	/���2 ���E�2���R��Cv�Nl�W���zv~�iF�	y��Y��n׏�E����LP����]IFGcI�]��za���H��yL���|��"����׋�+ ��i0��Ù`�aEo��Q�^`�'7�؄���'tLIɐ���-z��>X��J�Fu�]��.9u���Vᩩ��y�fq@ �C���<��~��򜅥�T��n��)�>ڦ��1 
�e��~AC[ۭ����O��J�g�k�;B�����G��:.���}�s�o{#a��gg8��C\5����zMS��������C�x���}��K34�MXykk��}s�v$��\������rB�22]��Ɯ�?F�}����G
qQ쮐��]��t��\\}m�E[�c|�㏁u�+o��r��(+�j��}�9�i� Qj��4�>��zk���$�u=Υ����o��U�]K��황X���|J#�3e��DpzKR���b��G����o����e�����?PE�^�c�*�x��G���i�n{[X0�]�w}yҌ�.sᛕ�0r����=gc;�N��;μ �эG��&~V/5�A�etqq�9���������)�d���O��/J��b�����i�\���������3����ᱠ�np���ݛ �����ʊ���c_������,n4�U5�3�k{���0%���u|�2�'�xÄ�/���������˶�P�NsXh�nf��GG���gMb�M}�á�{������C&S�M���������)q��-E�x�x�un���)�ʔ��}bxI4�����x2[o�<^0O� Pqz�������l,�s�˼099��v滶1��'��	9=�Z�G�ͪ�y/�}	���'�_x�����Bs	>q�mO
��L۾��YNr~�y�3:����$������Y��,�Ot	5l�	O 8�;53�[Z��^��������{��i�i�C��;�����.ARB@iiI���j��������ݏ�p-���������}�Y�� �@t�
��T;���6�:�\�c-��еaU��+>��d]��c����x�1�%*Q��.93T�n�S�-�Z�f~k�d�5�l���0֓y塎���:���>xmW�DJ�k�8?�� ��x*uKiY���-J.�����y�pQ$O�.�{�(z��8�1�ʁ�JM�IMs�O<��B�&8�Dy �R���᡺�6�׾��)��E�M��vU�+ZƊ�Ѐ�G
i>d�_k7���+��ը%��Ë��OӬ��א1���?C;L��w�+;�_k����>-���ZrC��#7��(��w{Ey�Α���:���x�gU����KL��U���5�'<���%Ixg܆���-���\�*�,G<�>��φk���̗�4ҙ�y���}�+P:�:hWwF({n ��P�!�!���E��?�n��=���x�y=�*�a����~��ҝ���[�wh9��v�6A]��:� !�|7�\<��y�QL�R2�˺ 8����Gy����-o��=�&ӚE5��ţ�s��[`9-��+�(�z�sr� Kt8;;3��wa�r�W��E>��ҮN_)��$�h &z;�FC֎���4@��U�����	y�kB�?t����cU���K�Gx8���Э�|�<Yj���s�6O����X>�lrrs㲵�5���7`RZY�&`���*\�	�\���e��Cc(��9��J���isG=::�ŀ�ORہ݆���Oh'����$^")���U��BZ�(�k1-j���z2��Vp�S���*�ݷ��\�~�I<�V---X.f��b�@�]���v
[��ns�7�1Ο�E�E���vU�����L��˽I�y���+b��gD��rm����
��Y.�	�hO�&h��@���������Yj�8��O3�EɊ��:k)L$��g���}Ȅ��,.-�27���~A��
H���J��b��u��@*��&B,j(x�@ wf(&������330�Kʲ�S��[�iN)�]�ƾgz(L�SvR�8����C"N��,&Po?a�)nS�}d��P)P���-�����W�����X� ��,�mCw�C����xxV	�^�IR�VnZ�Ӻ^�_�
9�r�oe���<J7�S�@_�~}8=_0�RG$�+�ta�\+��S4 ��E� ���k2*�;����e�1�3�Idw��AFb�*@*uuu������|E*�v X�S�_~TV��W�����"��o؞7��Y���@�љ|�jjT�?~��/�)��O�? ������e�Dqtfwww�7
/�$"�X���:�%RX�Ϲ�r������ߨ�o.�V�����2$:`Fl�J�n�$�k��_��&��Ȅ�4���f�fiߩ(}��֍�WcN,�bz �9�_�*:�h-�dp�w8�9g,kllq�_N�3�ck��/�U"L��V� h�p3�����Љ�l^?�!�\�1"#:��Zf�������P')�Џ\�pj�Ƭ>F����o�N��!�wP�ڽ=X���bY|Z��~�bnRPX��7��B(S�~�v��o{Lz|d�Ӌ�F�#Ugs_H�#V\̭P�J�:�@>�s��
F4��# ��Sޥ�hi}��.���b�
R5!��Ԓf��H3�����T.븭C^��H�� �I?k������ ��+,^�Ü�M�<j�p�u�}t@&d�Y@�#|��Rs��l��'�:dM�����,D��ɥm4���}Kyee/��H�<)���b�H�`p���g�E�:�3ps+D��ƕ��g�������nA���A6�b~�;̓�3���0�|��e�)���]���� �tc�99M8�U:�ʧ*��b��ZRQ���> �kY��E�b�����咶���5���T^^��ۦ��٪�	A	���4E@*f�߇"��0��WϤ�c�fr��������(����y�qe�B����F������o_���p���w��x
<\�DP���R&�Q����0!T���\��]��C��p;�Iw��A�Ug��c�����ݪ��o1ė,Y��pX{�D1=ȱ��Q���b
k��ϩ5?t�ӳ����e���7���D��{�KF~n5�8������r"s#+;�H;�O���Nÿ؅cj�<��+�~贂BVK_���҇
����\Vj�t����Z�iP���U�!h�F=J2����� ��M��� y��o�/qrr�[�-�1��^���*�W[���(��?r�3)��X��f'^�d�`$e�AJ\�_K� �A��������"sF_�r�Drss-k����oP���5h���	�#-���K�	z�����e�E=~���i^��nBy+��yx;�1>[���6D�4L�c/�������PB��0����_iy-��Z������{)u�����c	]߷�+ќZ������+�-�ɀn^v���I��k�����3ӵ�;dY �CHAq�y�/n����6�l~�����FF��Q���o�X��?L��;���w�%m�d�Or2��t7�j���"�������CLV ����ПB�g}DBME��3���L�++��h�IB� ��y���/�a���n��Mm�����A��c�%��~�����Ȃ=��ىM��^��~�
E�feU��ɛ��4"�1�\�]I\�*R�ջl�TR"<\N��y1�-h|q�}���x/=3�a䑐�j̀#?�����0�}9a.c�UC���x���c����d���G�B7���� ��=�J��)�@B��d���v6�\y@Y:��c�Ob�U����\o$��,�R�s'�00?�Xc�,h�pcc��nN�a��	����M@?�%��nϯm_^�c��΁�����c����y(9�v�gK��4�~�,z��3�V�xL�g�4Ɗ,���[�/լ����8ӆj�*q���t�t�,a���b�s�H��~-#��$BV����3 ���X�F���&��������%e���-��Λ*))9��-u94l�7�&fveszU���$�|+�xsj��Ǐ���B�t�����B �{�D�B4s6$�Kg����o��6��{F�G�"q��p�8��)�dF����5�Ym]��Ӕ��=a�r����w�q@u���T.($�i"q�Dl6��������M�=�z�z�D�w�8[2~��?(�����-
ő�`&v��x��E!�rӷ�$��z�ϗ��44_|M�I	E����C'�W��3d�uF
��4�8��|g@h�f��ܯ�$A dm�J4A5�>���;;���P�0������'�z���"�T�)%���&��ױCq\�bM����{/����@H�S)�3'�D�T��5����ɾ��l��ڟ.��'�)�)������J4Y�zĽ`$�/�XI*Xn5x���~���>̐�E� 7�c�8:�K}&�(FZF�-{u�ֵJsHkKA�gt���y� ���~ԉ��o�,A���TFZz��u�lG�#����x���3Ϳ$|-�����B�+)}k

�;q���fx��[�?ޫ��O�~�c�KuvD��K�>dK����8��%]k�/��4�I�K��]��Tl��ޑ��*e�*�v��^Y�9 {4��s6��~����l+(v<Z�����n,��{`B��{\�b���4��,��jI���fz�6;3ޒ���eِ��g�:�o��FP+��BW���$�!u�O$@6U��"e��@;5\Z�O�Un��ȸN���v�M������(UlYؤM���HTm-��uH���߼?z�P�>��r22E�ou�ۗ����d��ihh, ��b��F�$<�<�qd�WZ��˺?��ǐ�.��^�<lRA}22GF,�hs>�Ւ�VQ�k�J /���YZ�f"=*����H͋U��c-s�;��E��]K���ֲ�T"�3��tIXT��:e��U���WnM�-��lѴ�{�ê�5&�X�f�FO~ӠU[�W�tw�[f�F:o�J�K��z��b�[]͉Fk�"LU�njz����q6!��j�ÄջD����n}�f����l{��t�q�z��qJ��uXK�А�殯�5�±��TD��׮��FB�l,i�֖E��	\�+-�t�^����<;�ΜO�o�u~O�iķ'|μ�]�(�Rc��θц=��'ח�1+1�Ĳ\��Vuh�6�v��r4�a>�Bs_��B�]֧۶�ۆ�驫��B���N�I��G�0�b�kU�:�+"�Vo������y�ؠ���f%�P����l�R}""�M �^�e[���/�UX����VGX2�5���W���n���v���p&��SȪE�����k�H�;���6�@����;i#��x�Fw���2�.���K��o�ڻ����e�6�5�+�����S�-]֪Zd������3�@�������:�Bn��B�r��y�G�F�ݽʩ���^hdI|.��jTQR���tbJ�]�CcJ:���E����C�����VV�Nk�F�m��Y�y��a�@���B��T��������Y/�e\)�}��d���ѢBs����'n��Y��D?�������E�S5�u[��׍�r�!^j����)��^,�d��^���uʧؽ���}�aF*��,򵑥���$��k+��γ\��F�:����跓���Ι;��	�
+e���qv-�|�>"As�G�8��S�p��p"�|W��u���
 ���i��5��єUچ��@sA��ﶏւ��	��6����>�*��zD�֕W��^ �y� �,?H+I�Ni�f�Xx�y��Gr2X��Ĉw��4||��]����M�����c���uʦ���2������v1p��������'��t2��x���^_� �P�Q ��Z-2RR6�j�� ��N�K�����r��
�Ʌ�d�ƋaC{�S{��i /ZI�GJ��h7N�+Qz�5{�	N�s%�<�@�Ș��|�n�r��f`t���2���)8�$$=Uv�}��z�,���^��h���,?���T�R,	@ъL���S�-�����%J;<�����b"���9Jh���Y�l�V<ħ�#$��
��y-�/z+���H�M�ч�>^��I�|IDİ���'i0��t�����[[����y�`�q��.���gn��1ښ0=�{\9bm�#��.��mЇ�ߒ�ڰ(�������������=�	/s��Q0s�rݴf�"��B�Ņ�����pS�������	�Է>mMM$�,u/�E� ��h��+�����˰�w{��-�y]=8b1Qx
��::�x�l�nҸ>E �Y��Q����t��C�����ɼ����������56��@58ԡC6�%���bZ�JnM����^��ԫ��T���6	z�z*7h0��Q�����F�M���1�Ӄ��b[J����S]�BLJ=���5&/})Ah~R�L\�=y Ţ'�:~U�s�`=��'��π�r�oY�Z���]��V����'mPz��T���e�XR�K�B%���f�vŖ����ͦj�Q�dǝ���[����-�q����jJuJ-�/�gre��U�no��x&��*��g	���;bH��*x?�Z���{�rB����DE6�9�O����WX��O�˖���wT�0Ɍ��m���L�L�/��EӐ��az	�9]8Z���➔�x�Լ/���븜�����_�q��,�У <��j�^�J&Ӣ���W���hG[�]��������`.n|�|����u�jq�9d��ť�(Lȿ���j���mW���JEv����0��ggf�{��2�9L;�#�>�-����%�I/i����Yܲ?�׽H���͘�,�n�8k*+�?��N2���ME!���E���ċ�{�0a(E��~*��i��-,Dt�H2 3��¼��î��/Q�H^T�F�����v�x�s���h:P�P��eiӚ����f�N��K<� ������f1���}(=P��_;]6�^l��$S=j�k��{��<hqՅ�#LՂt��B1���b˙��㐷��rz>%6	'"*�w{Z��fqU���+�� d��Y���!�G�I�T-JƤ��3LqB}_��S�l�v�k�pG��2n I��C�f����#b�����cf����c��c�T-�Լ�:	~h!���]�Ջ��@|�<< �@v㛛�>��T�������8��n��R��Q����@��[����؞Ƅ��~�{�Rv�:���=w<\1���	11)Y��~��7 �����fѱ�e��xټ��&7:, ���ۨų����^_p�U��	���P9)�4iٹW#�CI��k֕L,�1~��nf����#�)���'L�%���������Y[~�%�"<���+N>��HdBy���Y۳������9ʀ�!�qՑȸ�~]�8z��"���K<��m>�({���LE�+$x�� ���li¯��w�rÉ-C�%"ܬ�|�>TÝ����;?�8@��nz(��<OnK+�w.�֞G�T�l4ky߀#�6���|�4o[�$p˔��b֌�B}��\�A������[ff�1(�7�\HMwwq�ӡ�� ��qG@Ȣ�w�z�̬�ut�u񒜜e�_K9]�Je�2��W1�1�����yj�G�;-R���Ű�?6�dH�b=7e�ʑq\L��e>�ֹ��?[p*2ϮR����s�������J�P������g�y�J����UM[{�1�J�T�А ר*�pFa�9ha!���Ơ<H԰��ئ�K�Faۃ��+?���A��\VJ��'���#�b��+�����g���P�`Z�8�Gѯ��7���$�*���1���S�n�S:K�c���v��P�P�S.�Xa�7�eamm~�T׸��U�v�]P�f=��z��� n8BO�m�?.�b8�n����hWMG��.V&3�֑�1��y�e7ӋJL��Ae+/��RF��Ɔ=�WWH�,F�>yL? 6͈�M�P��z�&�,�G@�ާT:�G�M������Z� N�W��bȠz?l�+�L�˧I���@:���K�B��E�����9��tY+R:�f�薿'�sjk1UE��TEo��1Q�m��G2jVέ�J�ee\p���zq�"�)��O�Ȑ}��Ed�¨��6C�A	3=���0���'�17?�P��җ<1)I�Q����O��1u��9���F���J?9�uJ	,--m멅��lmm�tX�%�{�5��P���wU��3��� ��.g����G�OSt���B^Cs�j�**�%���	V�������|6H��<��;�U�$C������G��t��`�4
�A��w~��<���FZ�����F�9W��X:_8Ya[��A���}�%E������f���x��-���� ��oϋ�����3Wi��vy�_���]���M�W�0�E9¬�.�m{u�)��n6�7Zg����0�f'N�r�����7�`>^n��=�V���B�vFә�_���)؉���v�� :��7���)��(Y��=���*����J�OU�����Xr��):2�Q+O+��b�F!A;6u�b�L��� I��vLi/�{-�6n�	��7l�`���>�67m�<C�\�gV�	(?i)�4��m��P)#�hX�S��z�Ƣ��'��C�g�Vo3))ħ�10��y���Y���������F�3@���Z���p����I��wB������`V4`��b���R��
�(��o�o���	��E�"L
RH7��m^��h� `~��a�� ��f�LՆ@��ݑsY(�S؂H`�e�xon�ޭm�R30�f6+ԣ�UW�2	��am9��P���;���_[v~�9�l,���xQ�lZ���6n~8�ps��$	$�]'۞mW3(D���j^M_��1��i�>&�����Ѿ�>�+�BU2�P��=�]%ك�=J7�>���xI"3;ỿ�%ڥ�[~\��WFOy[^�[����<�pέ��k��j�:�Z7�P�og�J+��ѧw�*��c�ᡣ�|���.�bơk��e+����9�!�=�*ֆ����m�35Ģ�xq���X��v�{����ۇ'QQQ�9 ��K*��W�.c�`�o))ee��4��<��gYf�Z�}|�z̰�#+��ɩ��Y�,W7Ut%��11��sg�Sww7�ߵ=��N˹��ЈY,�/��>�ԍ L�A!}?X�8�=;�
�P��Fb5�u�9�H��Й1+-P�3�{����]�|jz:!!�sL�J_��	�{��6���//omo�=?=j�SrZ��c�3-"3���R��n�X�����J
�� �L�tk�)�m����> �G����"89��`�� ���t�8���z>^���N�-��Ef?�\��!�э4���!q�'�|���F��sI;IG��ˡ�z�3q]D�Gq�w[�x��ӿh{�hO x�[�a���+�;0@+(H�&�l䪿����쯒��?2[�����4LL肙�*Eh5�1SS�qؘ��إc�JHK�!I ���|�O@��
�R	��������aƕ�������@�����mn^�lۖ�^!@l�^T�r�c2�]��˨_��~��UIhurө�H��?�:X�+���rq���[4��4)�_y�z��r��������HI]��*���Uqe%�5{����D��@��S7Uiq���i���!����8a�B�f/η?����r�m�!㴳����W,Z��p��eC9�d�!�L�	�ߩ�%������^�y��&cB[�DPf9�|�|�j��\�̈3k<R̼������s�h�Q���yX=JDi��A����1�w�#�.���&����^O@��[�N�/АP����oϷ�_�˃��_�x@�9���z�4AzS K�V2�&�M&��m9vF�]��G.O��͢���l����ѣ#��ݩw�I���Mj����a��PJK�Z ������$��ڧh�y�����'�8�'�-�KSM������p�\��� �l��>��miGi�V�sz�Z�;��5R���뾸� <�~qc��z���5B�o�4:�#�C{��)U��,���(�w�J�I�(�ex�d�w�K���`�kS�e�տ��^�����+ȳ��:3�@cZ+�tLO�T��4!�>b��g-�r��y�����g/=���9t�Dħ�lT'��@��m�d����@�}��zODEµ�X�譈ˑ�+�c^e�]��WY�p�x��~-p������h�(I��K���������ؖ�\����([fV.T6Cn��~��M}���,\�i��:Jr,�g�-�6c�� P�� ��k/���6i:�M�s*M��D��A��-��������Z}�M1"���k{���H4��������F�+�K���� 2�:QJ}C���>)ҟ��[r{ O�ntcd��;;문�����Am��-������is;��'��ɰ�2�Y��Mlb�K�>��� #�o#��VD���@9���)J^ D_�ۻ�$ (��o�6}����Hv��鑣�Ģ�N��O���&i~�d����E��"�����n�E��,��z���u@~�g㔊jN�޹j�h4�4�tJ!_�AQ�:"���W�⅊��f7��s�"Y˄���&��$c��e�-�p������J��b�@�/"���&x��g!��6���ΩT�6tD�/���%M��Z� ��
�g���G�t�ZX��),N�t}������\�O� M0�\�^�c9f������K��ځ�L"��7�~��Sќ����D	��%�F��7��z�ly�k��1���l�A�^C1�|Y�cIW��My|{��A_~39�NF������"ܛ�����7���2����w�n�ro �fq�ݼ'P��Y`u�3��<�
m��j"�k���s,�ߠn����nB:���~Zl�XeL=~"�N���Ӊ�'�Ӂ��]�������ga[�� ��۹:�U��p[���Ż\�Y���JD� �X�r�rl�r٪���W�4�:�����=�76c�ܹ/Uz��J����v�}�[��NFaA'8�7?��*mk7�2n�!�4Pt^��n.E� ee�
�^�;����TLo�����A���u�do�(U�P�cXOLx�S����%X&���)�$\�2���Z=5�t��9�p�.?�I��.�������;�~��ý�_�Ka,����:zٗu�AǗU���FlE�^��b��w�pd���%�0�,����~s��}FU ={5�<�]�6
��]'J�d�h()/G�D�f��_�d-�,8�9ی�MƘ�-|��z���z)��s����aɨL�7���漼�d�Oo����^ۧ�B��v1�Ӵ�`(�������u
o��g���ג�تb��B�9y<����b�y�H���LEwX�-־`f�����}o�XϚ�(��f#�JQ�x%Np�Z���# DE�>�a���G�Ov_w~��O@%�zDQw��ͫ�Z����8�-YS�S��_Tæ��)_Ս	�4d�6Z�J�$�#c9+-�߿s�k�ob��[���2��J���xQ\�����'q�=����4�TV2�_���k�Z���X���ē��OJ*�\�F���nn��D��V���K��7ׁ4��tQ5|�3�E�D��K����U廋EYJ��ka��1+�G����'�k��/�,����l[��>L�G�1
�B��M�����Wb�c�Vgtٴ^��~u���?1E�g� ��������`~�72��L�g~��/WM�z��"2Vΐ�b���*�B.��V}֛��B�N���t�a5����
�н\?�Vʜ=������Φ w7�h �Z���1{����vW�l��k�nG��,7~e߽۱���.W��:�k^�G��K����wGM3�W�|��]�c�^v���{=a
�'1]>@ ���IG-���H*|Ƕ�UP�o�1n����Ù��V�\�T��,�6PV�����+�_0���`M;�s��<�����trl�x7:u��a����E��b(���!uI�p��L�wgC�7�)11r�=~	����ya�m�L~z:�$�J�2��A`��{U���<m=�2�+��T�bA�!����$)���"$�:O�2��݅Y��p�v�V���݄�i��y��SJ���C^a�)��C A�n����TKA�c��'x�4��ZӀ�1e�r����a�Դn���{�j���癏O��!@c=9z�p��f��H������!��t�y��7:e2�K��/��'�U�������b���8�K/W�3X�<�~V�����͒������AhcL�J>���K��$F�g3��~����PW(���OG�q'2�Q��)NhȈ�:�̙������WD%0��}j��נ� "�'�zvj�?#�s/=�_�n�j=�0x�v!c,�w��C!����m���5��_�>.��Đ�:JP���7���,�A-d @!U���8���&%��ze���g@cd�3�?��H\�����5��+c_�6&�^�f~��s�cC��:1�$��	�p�M9m���b���B\0�q-ψ�O�¯�����xr���EC�Y,��V����;���!�	���9-�͆�v�zϙ�%ڍ������]ztr����]�/�RX-��>�H5���4Ѹ�� b�H���i�+�mWE��
��0��WfBd6�2>�n=]&8R!��(���W��_8t-AE��c��䣎�IKK[w�	�Ig�����"�'��G�$�����Ւ\X�^;@ˡ�s����\�:�S�_���v4���=	kbb.o��ɿU����R]O�h��S;=ϙ?l�_��vΩ�R?�pB��+����ľ��/j�cؖ�"�����'�⇳�5���9��P˲ݏ�b�=x*E\T�V��Y�d����M���F��~�wƚ�+s�n�	�eT[GϏ&U$-�g�T���~�AX�/M��ܵ	�b�� �m�`�_�&d�A�re��x����ϴE,���;�����> -s�9s[���p݃i���4�p�CwY�6�y���R�"onnq��8h[�m���3|���뉎f�ڃN�K@�n������ڼ@g�0X%���.���v憘\p�?�ެR�*!�x�Ɩ_��/r�q��ú3�C��Pā�54�P�)jz!���t:����hZj�J�Ԭ=���Ŀ������(��\��� ����&�ͭ�N�`|s߃�f�$�����y���r�wa�	6ʤ	�!i�U�n8�:S�X[��2�,nM����ީ��3b���=0k')،K�f6F(�.vD�\���(Fm�0&��Tf���l���cQ���X>J�
��PN������>���YD�(Ks)� ��8M��͈���tK��߄#�=A����m�u��؀z�ě뵋�t�qf�Ӛz�� �^e��S�U��ۇc������{~�ɪq��=��Y|W�C���yq(G3��5q�n���Ki�ym#�؂�(xu�o-ꟉO���#?d�z��Þ��"{�X��դ�d�>��m��-A��er��	C�fs�k~�0�%��X}��Pސ���{��Sg+���#{)����a�HS�v(���sM 2���]K~��������y|�����K׷	�>�k�7��_�ir��n�	��s���Eڥc�Hj��9�+B�&B��ů�/�_R	L2;V���U�c-��/��|��^)-qu���_��I���sr���)T
��A�[��^�IQ»�� ���M��u�]�#y�O�|�3�"чi�&�	�_�-���:�IEZ�:?�z�ty�G&��E�˩��]{��������?*�0b$��w���[#�Fq����S��oG?�e{�Ʌ����K򓮣6�WJ�=��y�\++"�s�4���h*���ȡT_d�c�H�m��(��ݭ�K}� �F�-� ��Wn��F��Œ�'B;!D1A����1�7��;�Ɂc��"�vDB��B\�c�MY2�fz���7)�L��q�-�+�'P
�X��z��ɰCw�P�̷c�Lv�jI�_M�1=�z���7AK�~.���a�A�x5vQ��pPYv�ӿ$y9HT�ϲ��u���D�$�f�P?��yp�
�2H�L��u<�`��k{��t�>�Vup�z�]��H���� ���@u�&H���.�;1����_��C�*��K^���d4�����y	$��D���H� ��������l�=��d����۰t+�C24���|�L�<�_�7ڻ��<���SV��AuTqvˉ�~�LlH�j_[������ �u� sq���c��U}Ľ��y��kCˈ˓��Y?D����EFYr�9�|�@9U��t0��� �g /��Y-df���y;NR-�o�Աako��#_��3�T^�V�"-��؈4�=�!MʎzI�oҖ["�=!<v"kJǡwk��oSnҖ����v�=�֪ϙD�c�莔����<�t����U����n�w�����%�l���]P� �z��q�g��d���6�bͷ��m,�����N�œ�~��4�u�a��@������ׄ���$��beZ�_^�{_��М���T|�������Cyz.Wh�_�~l(�/{�;
�!{a������Y��ޛ�Ğ�1���M.�
b�KwY��#x�c܎�j._��h��פͺ���ɲn{ƿRPF�)�_4�Tii~1^G�TkK�f&��6BL��,��C>��G����(YF	4�$�	����]�K�!K*t����ٙ���2�9���+�s��4ж��k���k��mܾ�,�q�Y61����v
KF�~9�!���5m<]v�@#���<e���*,��ms0���Ĵ�L��6���Ϡх��J���ʶ��)��
��u��S}u��5��S9��̂�!D�Z�t�ۆ�]����t���������F:���{Ʉ-�m��V��e�֨��8�nP�Å&l��*T�U[ݢP 	���x��˱���b�f���ذ���� �B�Ԍ�'�#M��Sh�4Ȑ1�xǹ֡���S�L��[	�.4*�}�̚y����
V�@��hƳ�P��w3*E���B�K���,�Q����k �\v��:�r}����ٹA~��CE���e>`����Ub[�3%�tJÀ�ǈp0���紙�IGB�;z#��p�ʌ����>���w	�Q�a^�����^R
B���{#E�9�O@(dՑ��l����R��9	M,3��=)T�&�#��ͥ��`
��p��{�t����1'���@�����i%��+�(����޼�_��ݬ� w;���݈�~�Ϻ�;|��ߋHWDs���*��'2_��x��@�4�+�6C��癩N������ �Ğ��s�G�^B#J:s�
"\�67�,��Q�\��B����#WD>�-pZT� ܼ/�-�����0+��(]̎;+6t�'o���+r����b:�B���q� ��]�T���
��ki�6��Y��Biq��p��޳e���!��C�ڤ����K�D���7`GD�F(���0�8�w�r��ފ�QbC` ��Y�����}VS$�;NGR�}��r��\�dVa��8���G���AK��n(6��L�"4����@ʠ�
�}�����"�.��^�֓AJ���&)����om~�r��~qb�o�ZS�Տ�3�þ���M��g��/�L�L�u���@� t耭g��Ƹ��n���ل���գ��R[i��c�Q�rk�
T�0�dj<�-�9�������'�H�טo5�Ԭwd�Y����S�!#�U�5�7+u͋�W!r�bȮXxz�|b�^�����>�����N�s{��9ϷO�����KSg���՝/����WT�e��(Y������z�=��=,��c�gh�B"v�_0�%G�����G��J`��	����]{��?&z!���'��������$8'����	S�����ZD��q�"I�vp6��Jo�^s{��_��[��ǲ+����T���Q��n�-��H�w+�y�y��������m@�`��$�ʮǱ��f�#�h?4`۵)gv�W��m��x҇8���Hr���Yz�s�^��c�p.�O��U��T��:fc�T����mۨ����Ku����OK:u�W�&M����g����]>���~1�Ϯø���O��E�֠�Z��U�?��m.+y�'�Ef����ڲQ_�z��,�wc�9d���eSq;e|w���yXɜ��v�|@c��)��i����q��b��`������Ds�I�픡ưq4�Tu\��7�0�nkf���=9��׫�(+>���6IIIw��ꓼ���|�sN�6�%ON��F״jc������옗d'T2��@�6EN|�+�J��qk{"pM�4d@�k��E�lm��HǷ������u��gO���|�e��A5���7`ෟq���D�~�~�/���I�w@�����`陠l�);D�n�����*d�R�����.Q�����Բ���Ϯ�#�M���a3k�^�&�3GX��:A>o�Mj�_@`�I�ݚt5L:O=�����^l'��>�'~���z���z��L�?Gym"�~'w�F�������,�ͻ��d��<��V�����ϒ4�(�3]�R$�ga���ӊr�F/&��wW�z�@�ɸ��������l����WF�Ҟ�(v�Yw������A�E�����|���̔���e�\19&6��o�.|�$1���qm���y���8Ux�Y��$����:��V�P�D����]@N�;�$�91_͗o��
ߟ�.�?~��-�·���U���4�����f�=_���1����fH��S�����Puu|�.,�%�pp�|@��W���1��g&�ɫb�h��⣻�>1�a�5_>϶����%l�|z�M�l�m�%�̰��x�%j��O��J8o��;���.-�xJ�U�����C�<ʝ)�z~�>��,IZ^�c�U�Vt�;����غ��z��MşG睴�P{����p�̋<>�>����W8Q��Koo�]��n�$�:r�T�?�Q���-��Uj�(}!�R� �,6S���P<A��Zǒ:����U$���/]��V�oJq_��ٞj�������y?@��}-���ęs�W��]�����9Ѯ����F˱+r��~u��������պ�����C�T��￥&/Ɵ�0��F��܃���p�G�(?h�Ѱ�>W�A��d��A��r���wVO᳅����r�?�-e^5��L�b��'P��,�iok0���4z�繲��|�_��6�����%����uptT��7�]��Ouo@�ɥt7�۞���uXrԔ����j1d?l1�U0��u�Ȭ��4o�0�.O� 6>��j�b:K�x������i��9�@�K�� ��Ò��QUO�����|��GC�1w�>zF���� H�B���%�Ӊ:�|Y��k"�棕4���cj��w����+��~���2^��۱�`�7I�NA�s�͏� �E��cW�gQ���7�=q�B��^6�?X�Z��w���?��;(���D�$�A�I2��$q�F%�!y�� �H�4���<�H�Yr��!Ð���m��>����U[Us�=�����t����no���%��TO��\��V+��4Ⱦ���ia��a<�v�`�c�q���\w�������]j�W�=圦P�(���۷��RW�0����~&Z��J�q�&�t�@�͓WW~gȬ�Lϣ���Y����hAo��%��Z��13�ѫ�]��1�'��U�g�����k�%�]}��I��@�n�"�A���{�:%M!�uﶪ|3g
AwM��B\�DsU��Ӏ��fr�n3>��c��I��64�������V�+�#��&�D�S+�?]L�l<t�[l�~%h���Z�I����.��5�:j���(R+ޢ�m�L�)���kQ���y`(D�-h��<��W.!�ZɆTO�o�k;�ް���r�1���(ƨ�Y�^ĭsR���\tbVK�Y2j_��h !�V�&ɀ&[�8���7i�'{d>c�y�N 5�������Ɂ xe(�����r�]Z�޽i��ŧ�T�����l5=/��9x
܃�wN�5�Uz���G�]�����Kt���=[Cf�%�^U�`�6����[�5m���u�|��#߶���ޏ%+mU��	j����Z L���R��UD\��L[��1j�ܴX�D�G��I��eg�0CQ�R�?��*��^%�_��4�|��"��s��QP}�FO����)��TAF�0��[ ��J���L~�諨*/ܾoAN�0�1�~}JL�t@Cu��s�y*�֭Q:kٙ���[	�j[�z��ߢ9�jk頟$E�;���ҳ�
iP{��^�CL�"7B�ܩ~�U���<��7���)��*���!41u"��q7*Qp�ۂiFc^ǎ�f��.X�F����G�|Fק�0�����6X�qK��%�2�tۦ��t~&X��5�}�N�&�Y��Df8������G1�t3�P�� �Y9����r�>�.ߊ}� |f��D���Zьa���0�Bf���?�6���|�1U+�0��b��-��gN?-/>����Kԫ��.�BF}��Ъ��"�ԧ��~��3U>��#]h�joyn���+x�9ժ|���TO��6Jm����u�y�v�Ww��g���D~!�o"t�LDv���u���Ԯ�N��`�NZ�눛X���(:aV��j�f���H�i�hd����ۮᜱZR�m&���Q��Cu�N��j]�_O�Zt��0��IL�A�og#���{r<:�9az��ae�$�oc�T�e�� W?�g]�T�������#�ظ�ޝ�{��x�Ta��bòF��C#D��cC��K���x�9h�C�%�%|�/��.f�ǂV$�)��V�����n������>{�A�YN��������Un�o@�ki`�Z�P�/ᇄ�{���Y*0vH���n�7@����2�����a�?�u�sHA=.R�ifB�ٍ%z��ck��xrۇ�3�O�JĿ ^ꌝi>��t֓�%���k
g&�ߕ�+��3��qؗ1�����{q)����_D�o5�$If��#jxI1Pɐ�o�n��/�փݰ��In��	��aI�n'�(^�]���
0�#|:�o�Bw�mk�����SN��?��ejKO�����WO\����?f�g�.]�wGg)X
�o�
ctqa��G�{�ش�4�}��K���.�E.����r������`�� ���u	���p�F �ϴ��e�;�����{�b��><ɒYԲ
}״����v��_Fz�&�s()m��Fp뱒Փ�|f�*(�R٢M�I�r��I �N�c&�H��bn�
0IId �W��W��wM���Ϸ�9�~F2	�q8�3��ov�;�L��DL�׷A�N} '�U��c6�Ǭ�����)��_g��>��X膘�s���[�Q�����ԟ���V�{���r+az@�"!��]ˮA���L��K��B��é���7�]w�+�Y:O����f{p��'&P���a�>,����w�ن��-��� #�Ԡ�]Q'�|�Q�/��Rt���Θ+lO��	�n����fuL�2�񳜉8��m9��nYJu�2�$�eWoQߺ	�����d��#� U���5��}��"�t�<���U����r�H���yj�|&��+{ +L�W���Y� ?�f;�����f3��Nkww|^���wd�B�^��I�� ��R���Е�{�h��_��c�v����0�TMא��e{G�,�O��SB�O���Q��:u����ዎغt�$k.���7�e�Zj޴%�	yW�qUM�jH5{��f��u|oY�ְ�+ġ��W<�������_�ɏVph�r����WG�U:	% �f_��Y�l� � Z�|�3��t	m�B����"Ԝ�
�*U.S��>�j"�HxV����BU�����~�)}pLk��N�tӜ���G*���UTT =�N/�026^�����4�Z��{K��E`�?zf�O���� ����?�[�Y��" (HfSyݎnF�"�
�$���pʋ���Ő;�k2�sa,�����%����(Ȧ���'�j�-�,����m&��P�����e��\&~�8
��pf�'L�/޾i���x��Rn!o��s�D]�y�'?���4���|cZ��k�UŁ�d�rg�Zt*�^�y��2��*�{e����[�2^����Ey"W�0O_�|�qS�Ԙ�ld�3]Ű��������vZ�Z�sH�}l�� ��Nb�����#�����+K��jǩ�`*� Q4�/���\��}�1�T�������Z��I��8��cZ�~��.3���43��Yx|7*!5�A)��,	��B,��H�@�u���s�y�˪N�7[��	f>'��͓2�ٶG찧��Uÿ�o,G���8���s(�b��j~�bT�ZC.Q)�Qu�D�ߋ፛��3���{�2��`l�>�Y�j* *D���M�t�;��̄���^d
%j�$P �6��WسŌ�܈�m��YR	�Ǉ8�
�'�*���6�2�P��;��O�JZ��G�ɻKw�EV���D��:?�{���4�z40�R'v��g�8���d���G!���2-A�)��)�䪃.�i�8l'KYiE�]d�����p.�)��+�����-�X3�Av�����^���^auF�WI%U������:Hz��f����"�\��'*,kh�	�9���$V�
O�MW�T�	��v:\$�`<���=�:v�m����u�榅@��!������u�n��XˤrN�xKvj�N��1��0�V2Q
ê��
.�k*Qk�.�W��@jw]i(R`�xV�)ϯb�Q&���_��N|�;��`�9Y_�E�c+��?]����Y$*{6�oޔp}�����%+�A%�T{�PY����q���(���Ӈ�#{-�6 ���6Ocvέ����
T�M�E���t��y�I	�]�?�����v�7`������z&(�W�Zx�	"j���|���۷}>A���vW��s��ͱ5R?�[��$�p��^��O X�+��u�LL�H��g����p�ɀ��@<A=���4�����B7W���L��Yl�F�[�R����9��}�k��5j�f���7B�JG�AZMN�ȧ#��8k���Q����w,O"O����?���?S�� #�*Z71�HɂH�솽΁b	<�}&���@�d8�:��eQ����˴�I��U#_��H.U����LC�i�O)�	҈�ȭe�,�s�^E��ڋ'~��y�143�����u3�>f�Ѓ��h�ҭ!9���J�j����?2��sT�� ݚ���s�6��#uG��$��$a���̫�?a���\?��$W��7�ʗ�VB����J��%aWoW��A�V�?R�7�I3���j
xN6LM��+10 ��Ql��LԠ��<8qq-����\�1���sGG��Je|�d�yeڿ3/�_�����[�>��#l5z�P��Ԥ�֬����ݭ�\*���Ϛ�@y�8�����8K�D(������A\R�-{�0��G�?W�q	���fԂ*d1�Ⱥ�ټ�Flo�X��C�c}e��~��G�y Ӝ�铔��t�ƹ%O��[6=�<�J���Oy�)�O6�e̟�ǧfs��r��O�bxdKW'7�./�s�ˠ�uɌ��{���<���*풵+��}��(@�B��'3ZQC�p�2d�J��JһEP��O?zlOS��T�As��������+��:����L�����hq$_�YC�X�Q;�/~sj����Z����!]|��dqa�Mb ��o�@��R�K�c_kJ7�t�yc�dA���׆P1�o|*[�~tl��lCy��|=L2���~Գk�\�Z"Y:Gϔ\���q�.M&>���2^dC��'v?5p�|4�b��^�PY��|~G〙�����3��0Ir0~7��H~)t�^&�el�j{g�RZ
zVK��I���E[T�d�{�d]�
��P�U�;��x~��?�:G}���8�D#@��-�ӗ�Lq�o�#�}�G󬵠��-�y��]_JhB6S�xѹG�"�n�K�a/�ǅca�?�C�9�T*XOr	�{�vߤWaUE�M�Fz��a�+t.�����qɀ.׶K���'u�{�P�������Y�$�M�~&w���QR~Hɦ����mF{_�ý�� ��㝭���d
B�m��+�=ZS��Mb��I����Te��]O����*���[���B���8�Ql��R��ψ��5�o~^mf5�#x��u}��sB���3^�^�����T�`_���F�U T^�wy�rW�˥K�y�Р����S�g}���~����`
QS��@"Q6.�8��.��0;� ���7��k�B�uh�p��+ǡ{��)Q�ʽh�*,�L���^d���wƹ7Wuid02\:�xX΀J�. ��&����X�T,O<0W��~�5��Qi%o�HQ�%/�����&~�I�)������P2WJ?��P��d�4�=_�l@ ����er�,���sB�v��	��;:�"S�쳎����t��-^�(Խ>;Ɇ2��G^�w5v�Y���h�3ezs�>^�Qߴ��Z�� ���H�w6����Y�<�
[h�KN�߭��������Q�fx�oPu8�"��RbFp�s�� T$�]~����Uˎ��,I�)�//Տ�,U����� �S���u�K"/E�xnR���	Uh&f��h���oVa��S^[|c*Jׯo�g�6��Me�)���C�) ��b��qf�K>ݢQ~A�t?t�K6>�u�[����`��2}��U�ο�x�����u����>@������^>�;�!x�1t�+��y��ً�ȈZqތ4c����;
�Y�o}Ȉ4o����F'� �>�N�&��NZ|#��
Q���F��e�%%t��]�~x2���C��<
� ,��9/�\�о<FHT+G��g�s�����M�M��M]|�l1>�o��K����n�R�Fq��X�}M��^E�fm��v����!��O�@Dx�'t�������ZO�ӟ�J���f�u�GU�z3]�7`�)#�06x���j����`�`j�[9y����]l�DłmeuBS�Ѱ��Yԭ����T�:G'i:.c9zS��s� ��dhV�P�r�%�čX�{hH���w
kn\zC\�[�H5m�a��Oiwk��U�}�|�7����}0���ݰ�E�1��r��GUݱy��<���m�+��ʫ���o�C�$�⪢����s��/�
�+7�Yb]�'yX�'��ҳ�}�T���?��|{H�����eG�2J�e�S��w�=�g3tۜ��テ�v�T�9^� �jU�ͪut1-��Q���ژ%d�m������b�_��F��!O��4r�X���6�`9�&R���C7L���o&�,7�`�9�f���w�5n�ϒC����+��[%����k<����@����4�9�''�	��8Y�ɕ[_���3�c,�I	�% �Ԭ�B��T4�)?~�׿l9��E��I����uȈ����jJ�y���ӎo�����_f|�v���RP�S�ii�����I�ճ�/��*��8�86����e�������H.�>I,��sy�͑��h-�8�x=�z=���IK(al>?I2��D��	�e�`�7�M�iZK�rԴN���Pf�֧.�m����h���9ި�k��f%wԮ�1<�
ww�ˮd�y���4�ē����p��u����Y��"|ٍN>��Ds5UbC�i1��33ֿ�����_�h!�S֖0J�b�Q�|�e�����|r0��_?�@��8r_�0%/=<L>ޞr~�^y�F�K��:�(�'�����?unf��{�g����.F9rg�"
�`:v!��*B]C�&L�p�r����'	fS�q.@�24�'�6Mr!v�Hsᴯ�y�����fxw��-s4����5�I���|լ1���}�{D/���&-���4J�Iϳ`9�f�z���	j��ox0JЁ�i>��8D�c��ǵ�!�: �]n��B�Nf�=�^�N�%�:2�u��}�4u�y(�*X2	,�,��h�Dy2� >�[\[��'/��U�̾:�Nl9�<m��%�nvh�7x�w�ɹ�z ��f�V��A���kf����M@���zRl}���)\q�P�=���c�VS�O��1>O���΀�`ӄ�l��~Sn}���:��%N����_��\�T���GtI���Ȑ�i�u�c��9�l/��=��w������p�)@�������Z��U��qѾKd����GX�DM�6t"B�!(*�wL��J@�(F�k��ŉ$��=0�f��-�}d>�Q`�W���YP��y�Hm��G��ğpߜL��E�Þ	�bAHu��M %��8U��MG�0]��Ä$�ϩ����k7�|����V�II�Qж,4j||ąs.��7O�_c����|{�n�N�S�����3����M�f3�;M��;�3�sP��|6Q�8��m,�b���
�����ሰ{�_��wQ؃����P+�c�#�ыL�{�U�-)��Nuޖ!Pq}�+��/3�{�{��6k�3�߃�?c��ǋ;`�mYm���UiC�{�׊�_�V�hi���7��
�p�8�A����Gzy�="�qӤ��MU*�oy�\����]��mX�;�����@>����A|H@T��?�?�v[�Zy�%�n1��Ylk���߹9�l�՘r@���Kt@ ͧj���nN^��?�����o4zy
�u�,(M"���+�x4�(T����]Dļ��L���96<XMM���+��zuՍZ
Ro�h�&ז�"� �317��E��@��a�5W��B�|mE��AN�d��,��.�
Z�*%�H�]��O;^9�YSA�t�_���B�:��V ��А�+�w�a ��DY-�n�7���d�L`ơ�GXW����j�N�%>s���\�n>��\�a���JG �v�d*yJ��j��b�L#Yi``��@�RV�+�T���	�7�+���@��v��x�o���M/�u6f��5 r�ԵB����f��y��Bep�࿳��'�}>�*#ñu'���,�=����!P`����1_0l��[� �_�L��&��^�H�h3ʉgb���j��4l=ւ���8}
��1XC�T��;���Ֆ7��dԛz�=�WQy�K��6�����y�z�
�.��
7k���
�$��	����+��������5I4㳥�X*�WUy~Z;�n0|�	Ҟc�����Rg��Z��k�e%v�Uq�pG�C�B������ޮ��=��Y�����hQFY�B۰����Ag��؋�K��Q�Ȱ���5%hc𫶹�z�v.�<��ޏ�?���哾��,J[`��b9-uW����	}����*���Lېw�)��L���b�V�.mc����s���[����96�-߾)��� -Q0*�8>浿Y�.�@��ܼ�}��X<�e]��4Ԃ*�u|�GKV�l��΂
|�4�;�3����Ib�sf���.z�����:��m�x\��`�6�o5�󱎳ɫ�g�y�E�H�ɵV��ȸ��RA�T��z�ـ^���5��fr����tp�8j&?��0XH~�:�����@��8�9Uӳ{�%��m1��>6-���W*��̲2�J�@��Q�榖��g`$�t���Rtj�b�S\�	��i�t�|��1�&2������?��`����}6�	u��뮜P��/��m̓��e�l�aWi�-��{��Ѥ�C�ga�����5,�8�m�Z�Θ3g�����W�s�(�U�`5��Xwg�@r�PԖ尔��wPA�8Vo�HK�~	�;N�%���OA>��vo�C����������c��?��c��}�w��l�i$�|��v�ič+Mմ�"��?k>�?���*����W:r����BS�q�V��j��wL_�*� �I�p������E�ys�o���}6�&����^S����0<E ���~C�4'�LrҕNb2�	B^��r&�n|K��Н�Yz:��*橗�KC�-���'��0]�{gI�x��*�@Q�>T���?r��r���fC���6&��C�r��v3�W*_Q}��ε��k��o��� �q2ҥ�Z��]�؃�0n�6�>��|7��7��0ߺEOb���=4�4#mp	��Y�<M�1��eͦ��K�~�Eܨd��������u�j�(L�>�a�T�`N��:H8���vm�~HT�C�����|���@�qJm����>*��=�jY��4d�:�hh���T���7>V�O&��^z�&�v�}>�|�=���kP��ډ�Yi�]��m�*x����6��j�|���h�Ӄ6lu}�ħg*ŭ���5eq7�n}}�yʫ
,#o6'wMy5.�rV��xTGm�(�b9��ݱ����� UJ��$� �D�䄝�򁛷?]U�N.q{�3�`�ț���A��ln�T�3m$*�ӐĽ��Ԋ���a���ДO*��8^��xH0����	1�3��є�c�y��C��˭��C�W_�nW�٩{(��{$,y{�j^���h�u]!���sX�V_�SV�Y.[?{S�gOW��
�o�<�\��}�U�ba�&�S2��Qe�"�d>�F,J�.��I����nh#��(����o8Q;}�;k}v��a�scXP�#q�cp�B&a-U�Y�D'�l�gY����d��7~^v����씣tϽ�ߋi|�r��3�j{�MBy�	�����W
�xnѩN��e�:�ᘽ?�p�$�W���M�	[�"$��3꽪+�K�m�Y�W|J�ben1���{N���}d�&�[�ͦĹ���-X���e���2!yR�'u�?NW7�4P߃
�x���x;R\���tԠ�M�s�L���h�v�۽�t'd��;�D�R�����Vhn��<���	2ސrou�	6�� �[�&��Ҏį;	�gM��q*t�F���]�.,0�ͽ�_���u�����ѓ�/�mx[��󔚊��+�*,�FP�Z�S9�� �S�.C�;�a�s�����׾���峷�~W�������yv�������n�m������TQ�+���fgp���)�;q8�~�r������1�/#�N�K,H��PvV'��b��Iu���Z�Ӿ,ȴ�X]�~o�]�i�#��f��}L
�="5r�����ɾ	T.��i�3�k�������ee]Ly��8��s�<Ĩ�"�@x67���|�&t��e�w°��Q���%AH �^��,�\I�����f��ՀNM�K�W��r�������|���,E}�O%����IqUT�!��1/�
�#�^�
La��P)_"�4&[jč��޵\���������9��90�A���g��3��@��}�)��;�w��!����j0�8�k*�Ũ[꒡O<�;$7�_��t��I�i� �Z��T��X���V�k�C���=j��~f+�3;͢ ����,ϣp��Ad���2���"�8�aX��\�07��E6�`��@�s{L��F_{�d�X��B�1�|"Q,���M�f���@X�������_������5:�;�(�$h+�n����`�^j��!�a�+��ŅX�{?��A����������ϲ�������pu	$�u�N9�;�*���(K2c7��}�ʗ��`�Y�f����+c\��ω�>�؊Ԙ����}�YY64wIW����R(%n��Z�h�,AM�]���"-�=fo&���aoǆc�}�`;��B�?-�!)Uhىr�+�vG>�5���$e���^��"_{�O^r\eߩd|a��$J\|c��#��Y|�~��i���<e��*g*A��'<r�0Z=Eдk�r��H��H�cK��u.<�������Qʟ����dF�X�(���N�W�֘5�� n��������G5��Jeښ>S�1��N�擙�jE%��f��t���x�!�{�Je��>Ԗ=ut���e����=�P��Q�ŏ�r��z7Ƭs����gD��e1A{U�p���wڟ��ز�L�F�f�I��l��0��g��(DsZ�������O>N�-Y��u��w�?�m�N��uV���5ƄԴ�md����ݛ��g��3�i� r���V����4�R�~��nvn^7a.:B&�_ʖ?�e����G�S��S�hm@��5^��`�?��Gh&�zz�ɭ��1�e�����B&ſ�,�����]�^r3�?	\B&q�FywNҡ�{/c���pd�hޭ�_�h�dJ�V6���b�כo��i.�F���,�c{�eG��ψ��{�\ �]B�G���Y)}H{��	�Ż�*s��u1���s�\�ZC���q�ǋ�OJ� 0���D�!���7�� �;*�� o:�R�w��.�N�e�����.yQ��rCŬ���1��gcT]���j��>-�0rOeю���G�~����>�ȗ/���3�
1�R�P?LE\ ��ܴzގS�K;f|`L����:7�d��q;�@�}��]����H����X���o�oD���~̺��x�l�ݟNb���}�@j�S�:ݒ��lv?gs��g�fr�vXמt#<,���g�'OD��`~��/s�����$J�^�&�'����y:	>f2����SPI�����% !;w/�A���{�5x�%����^�F��h�9�NÁ�~%�����n�T�����%��>IKض������m��Un�E��h���}:�?z�g�6�4�����~G��C��+�k����ǣ�Q�n�$�w���m�1FF���a��u��J�;������������ɦMhe���Ԍ�!,z���6��F�i�sQ�=��i2Z�A�K����ñ��	�@�6�����T�y��9<U����@���ay�wCs�K��t�gh��L&�v�LZ�%�L�����(_�(,c��!�^\�Ñ�rndU2G]v��-D	U�7{�%�2�7�� ���p�"��o�u���9-憎;�<�]���s�7�Ӆ�,N� ������8I}b<;�,�e���<��i�ö[[ �alI��e���ܞߜ`����\8U[,���{�\����{�g�6�?΂]���ѓ5Ż;$�����Y�Y��\Ue�~���4�~�1�võ%�#`����Y
��:�&�~)޿Y"�;��}~��U��h�gu���PK�`;�����!��n�6젙���Ƶ��
{�����ˬ���I_Q��+�_ !k��,��0��e�Yi��a��Y�u��������М�a�+fy��b$8�8��+R�8O,�G%�K�i���/PEg�����GcoN#d[�O�]9>�~G=$ƃ��\�	��|e�����M�O#Vu{��xR��~���!���6�s<לO�w����F7��PN���+��D��wO��ѥ<���)6�ק�ţ����I��7m�+�:�G�2���<_����L4�n�b���Ň�@�B�R�PFF��B���F��`1k6z���;n��R��W{���zc-K��g���\�/.�k���b[0R��h�u|�L��Z�W����S�[��1w�l��'���K�����#�l�d�*!�8Ze>{=/S_�� y[����t"��P}�����U�?I˪Pp��]Pj����Զ�dZR��̩}��~,=�!Q���h@��A�x��Q��d����I�3]F�}���E��p��|�;���ix�IJ��h O�ƥp�D�fP�q)1.�S݊���|�Ad4�ڌ�b�o���� �n���_��@/[K?�4���O>	~����	�K���H7�*�C�$�����y:1jn�����x�o}5��.��B�K8۰4�C0���h�6���}g��B?����%b��3x��z�+�%��(���/�쟵���ܯL�2!G�jڻ�N�f�\��n-�u���y��X�ثC����I�5Ʊ��a�|�_���0�_0!K�ڜ�~�fF��tj�F���/���̀�2��-�nZ��ݰ����v^�df������#�+�g�	�Z�͈�U�m]F��w?�!R����!��o[ i�^L�	�r��B�/X�R~�Ȧ�/����	I�$��i��"E3*�#��d]��Q�����ggg~w���cb���G�Z� �[�_z���'��8��"y���*e2]��:������y}���黤l���(���+�|��Ds�"�K3omO�	�Z�k�'�쵓D-�I��b����%Ļ���F߈�Rw�ٿ$�,su��gG`���뿋��!E��8ݻ�2�T�I�9?�ا1U�v�X����&�+3Y���+�W,>��')j��v��"�E'�EO�pV,;O���t.�f))v%�! �(|l��j�
�ؽ��4Fh�pc{$��q��gS��ݚ��i{Kx8�ej*ޗn��6�:��,��V�M�`z��^��
M��6h�N5�V]���a:O{�M�d\��ީ�w���ƬW�g����-���M:]��J��A`5o�;q�;qг������Myf��e/-�q�K	}����[?�[���	����Hl���� �ʳgR�Rn�e<N7ȫ�z-�9�bak�r6�;&�r���W�n?WT_x�0kPoH�����Y ?�]3v/0�v!���6-�RG�����{�6�l�"	���v��G��R��Hg��IX�{>v�@���F:{j8 ��;���������i\��y���C'����'eˋ��맙�>ȩ����,��M"�=F��Y��A���LY���13�����P����ݪ�[>���#N�D�x� %�'�i~w��I�p�͚rf� ��)�1+Ic������]Z�/:��wM��W��""��Ҍ\.-�.Z9��@��RY/�>��mh��㨖�J'\صyZ�o1���Z]O�O��~�H� E�@�x�Zs����{�<��ѿ�j��.�.��W�M�n���7.�?��x)]����oG��$��=��[|T8���{�{.��5K=��{�'�z-;[����#l�1"$�J�G�Y�qk4��������d]�k5�ζD�^Gvw׃�(���G�����������z�S���f�~>b�ѧ�fߘ_���QK�<�y<�Ѕ
azC���2��<Z.��0/�%�{��Ki����n�7�j��RE�O��.U��/�~�� ���{����F�3���ל��ɣW����a%�;�,���<$�ck|�|q��g���AD,�����sED���4�0Y��Q�P}��:��%)��q�|#������y�o��(�}�i.t��60)ߟ8��	�طa���^����U��Iz 	�+�_��iH)�G��ߚݾ� �Ө{Y^�OZ�WD�^	��?敞��>@�l>�Up��/��[��oPk���~r���A�z�`�Jhԃ�~��If)�h���x�J�����k&��s+:�Z�kj7����L�'U�Y���ͰZ�'�������i�J��ly�(�{�lr+���w�Mex7$T1&��W4,oU���I���<,��$�8�aͶ�$	 ճ)nG�{����c[�;9�Vz�$*�w��o&&F�b�~9vj�rM�LJy���GKy$���g?�^���LE���V"ǋ����9�H�~�J��@�u�~��0���!��m�10\���q�l}���0O�*B��Q�^ �Bz}�̘;Q��y��f�^?���Y�>�%��`+���mqw���K�={��_F�܈^�`	�������=ߋ7}tk$\���h��8z�D��>X�_4T�՚����q¾�~����k�o��
O��#��M�Z����^/���Kq{1I�=���^�pa�E�CR,�`�߁A�)rqc���㤪�A��u���/����U"�[����ޙr����|��{T% ��/�g���i	}DkD� y��qg���Z����|ז&��:��>�H�W���Y�O�MV��MM��b�'��O�M�̤��D���C_�lmʞǅ'�(�ƅ��D�E$�CSQ*����^::G������My�K��[u��f���'�Ψ�8J�c0��;�޵H��L=������Y+**r� $%vtOD؝�������4���u|���|<?^�:��F/w��j߹����A}��=�W��>�h)�[��d�����ۈ$L��'[�/O�^�쵟l�8�om�ז5�tbWA����V��{����z���GZn�{3l�x;M�k���$������bQ;���_����M�¢�������I�w:����!�i��sb�Z���	�P+���3�����z��m'W/�xY��I9�G�-$F���5��B����}.��wKX&�O�kfYX6�M�� 3�c���\�r�٠}���؅�7M;�4qG���a-��� �a�ֿ�,�o�5\���q��}��U,��W�>�߁O���Tf�N�����B0��s��ƹ}ak�H�S%Q����spݾ�s�6��6EB�V��~T���e�p[�2S��_�������Qj8Ϟ���1��b��`%�Cgo%�q��d��t�A�5z���h�`O3���&ׇ�G�.7�w�B�N4tU�8[/�t���A/�ɷs@����_((��p����;��#�f?/+� ����_Ӆ��r%ђ�g��.��������[~���ss�bW�d'�=�¹�m�ur�]YG�K��SK%9�X��|���n9�W�Ƀ���QM����R���R��8��
?�Z%ɭ�^s������?��)�bN���l��b���蕱;j0���݃�%������������Z�Szi-��%�J����=�}��keZ"�������\�K}��F�־��qa����A@_wM��"Od����`g��~�?V�Kz���j塙/ث՚��^t/y� �d8��$��k�,�ձ�y^���op��-�h�Ud�enw苫���P�вj�"�����I��W)�~)�9����y��V�4e�Mnl������t=�%�"�����t���-�}�R
h��&��'sI�?�k��K!2�S{��O��^3�`ӹHn�H�:{,�b2����P3i��\�8c&ԊN4�|�k|W�\�h:�:j�%9y�#��`7���Z&�M�5" �Ƀ���Z���C���I�Y��k����|�r|��P�(����쌓`�|��3�:"��]j�O�%���ۊ�V��v>$U��D�`k����e���bލ�/��9.xR�fu��_�,��*F�D�p��~n�x������d$�}��޵~�d�q"O��v4���m�ga�g���6r/9��7k:�5=LtعM���T�`�����i\컸Vni)߼�{�9���n��l!8�F�/�Y�C���Һ6����	�2Ȇ�K����O@,[�I�3�GW��A�v��T֡��\	0��=>�h;�����Rҁ���+D�/nw�����4����jЅ}w%���tӧtÜm2��=򖚺����^�b%$�L�Bz^�SX��O�l��w����O��42�C�XZJ@ZJ$��Kx,�H��Rt,;�2���3�@T�_�`o"�jn�a�;c�� :�V��ysk�'��d��+M����x�����6������q��e�z܍���Jҝ �0��t�ߐLs�M� �Z�߄^��/DEo����%�@�l�A~|����z�}���)%�'ao9�{K�������r#S���O=D���n1�bk��s��������Gϥ��T�SƆJ����lk�:�����-6'k�� u9c����{�k]�C���<����o�uZ��C�<B4\�� ��^��Tn��~l���[�$hA��[��k��O�c�W ����wM���5ɨX>����*���8D��hq1����̴�ƻ�&G�\F睲'f�,���W�ө�	��j��f�ÿ;�# �1��%�7�~�Dh��T����WƟ����#-���o����X���ȋ$i�'��)�ݪ�	�9u4�|Qs�$$���1�Ѐ;8Z3��p`txz?�!���TW���ǿ���D���"�(� �J߿�-�����"�G�`;Y>��E��4�������w�qj]�r��lR4�Z����������_��]ca�:&�k��!����\���0��ږ���G�\�.d��wH�X>@���2(�&�.�{����n	�����<�{pw� �!آy���U���?[s{�{�i�魻8�;:�q���Wz��ZE	�S�{m!U�ݒ0T���.�JWg�N̾���l���ZTs�B�S�|�b 90@�|�o�Ny(m�W#y���u���!TX�u���{M�#3Ӣ�ۉ��m,�	�;vE�yG�h�8~�~�Hj{�[.��H"y:�jĥ�գ*ޭy�g�B6�oI0`�
:�y/<X�	�}ݬh%{T�z����j�<'��>,�Đ�[]��mr��!�LeR���G�[~	3"q���-A^�v�̀g;�@��D���_��?��>~߷;��O�R��~���L����#	LS�(HA�G>M]S���7f.g���	��ri�p��g�=���S^Ə�D�{I�6h�6���W�9M�O�u�+d��,W�G��t��;�Ð�Ϟd#���v�
}5�P��%��p�qL��ۤZ�"�5���W�B°|ZT-��z��D�B���_��uWq�Ҙ@�x�5�j�+�m:�G"�� ��r��L*�r觿yV�A��$	�2|W=�-4w��
�}�Ӧ ���L�Y�NMቷ���_y�E�����j0=�,�O[� J�G*T����f,}tUmћ�)��q&N��W;y�{�Q~�kGx#�ҙ�մbj�-o� ��:oW���˚`�P�ö*�sH-�����Ą��%@��?2[���D��_��H�w�T���B��+KI����
�����o`��ޘ�>07�By��I�7n�ΐ2��L�#Uގ-���l��}�o�}Y}�"�����^�2�&2N�b��9ug $�o!z��l�����2Z�z��}(���u�:��%ڀ,�ʒ.-l~�AX�C2s�&_s���U���թ������'ɲ=J���6w7l���+\��D�	�zќ	�Dspk�8R;�)0��^��_'�!�n���!g����?Ȏ���	z��sx��q>�����;��^�5a,�˝�r�M��|�O.��\i���F�f������>���������䵋�~�&������`V!�����[��~��n$Xwނ�r��;���Q���}�C��Kp��$����@�׌��M����]�g����ex�m)J�n//)���ְ��q�����G_�f�a�t�wꢈ�Z�z�#V�n:�H�ݿ�qE��vT�	��Q�c?{��r��dE����!�W��1��Ls�ş�A�����˰� ����ۻ��^�:6��_�F�I�A��hzȴ_���t*>2�%�7!q<��t��1����1XL��f�:��vA�@e���X�	���>ڧ�˾��r�����Â�Djt��HӺm�7��[��~P㗗�"�t��b􅹘`��xS��v�O����h:����� s���yz(��Q����M2d�_ l�-7),�{��	v��4"�dײ��J�񖞛}5�x���z�C����!Ӣ���e�*b�*��(��u��-���L}$!!��<��
���?R�3Q��C��W%�;�J�"u(CQ�g�2đJ�ɻ`���r�]e�l�!5�i�������?�--,D$Ȅq���:�H�A^C�on�� � �w���4/E��C��{sf��(p��
�u%l�;4�t�uBڕmx�v$���Qb���p*e�i���p�	�[�����k�@�d�;0Fp9o��5�|d}�����<����5�@8 �����ܟ��Q^�/���8��)�eǂ�x�ز�l�Ftj�Kt����+�����\�m�fJjrΡ\�Rl��Rf�L�{���(M�E5��eE`�{��0�w�-$��W�>��7B!��C��J�������n>��;ګ��//�|G��?�$]q/ۙ���Z���۾E��zE�vk_��A�MҾu����!!�D���Y�� 7Kx<W�����h�n�8��Y(
یH��U��3����-ɉ�PV�U���\���m�vQp�2��!)�n���������/=�D� i���H]'�=��::��q���aDu�{2�a˓%�1��.�]������!�Ra�ǁ`���Xf=Xg��HX�����QށST�}�%�&,-URv �R�©�	�[=KQ[�;�J#�.L���G$��MB�S��T�����YJ��t����������]n?��If�m���k$θ�6ɲl8�FW�CcA/EW�
!�5-~�DЎ�5}z+�WRr��>��`G�1�#��;+n��κ.���$C�*5J�U�p�j7�s6��}�xHqv�F(KD��d/E�蕹 � a�_�갶څ�z���|����]��Mơ�+l8��p��e"h\e_�Gs�*���Y�&���dF���r��%s䉲�߸�W21�9���}
�`~���b^F�3�5H(�D���� ;r�mߢ�˦��j��ߢ��{�Fl�l��r�LR�g�R3΂�3A2�j,T0�b�Jc�z��Z��i�ãۇ���l�COSńp�R�uIa�?Q_��A�����#qh2֣:a����@Vz�����z|&+�2	��[S\��3\����Q�p�g�q9��`?��.�&-����/Θ�B�qF	�F�|Q#�a�OJb�ðI�X�A��)� �|����9z�#�z�[Lt^m�u9���J�gR�YA
�*�z�F����a_��[a���g�}����ד�_�7���߫Yɬ�;�=�!2�&�C�&J�s�%M|�G*�ŭt��~�M<GqD������UT�uj��w������6ǶJk/��E�����-�w��N���V��[s��"�c��q%��`_�J�|�+8ǟn}���k��Y����&�a~���Ri��/���ʕ�n�K�:Ip~eK\����$K��]*Ȁ|HĪ'��ի,�2{�ƥjݻ#���\�|\T/�܍��l�Ý�@����_C�i�%=p
�Dq/�n&���*_�U�` �?,�b��Ĥ�1�MwK� ��Փ=su tTd�悴�-��c!3x��H��yu�T;i���Y�hj�8�
%u���i�P�� �yS��}���Y�����<+����P��
�+�����'�r�>[��
O�U�� ��5p�E�s�p��-��)�g+�#��j�7�CѢ�C��h�$Y	7��AS'<�L��F�����Ϋ�%NA�d�1�'�\������D^{��������֦�q�支+��
z�e?/�9����8�� /x�\��j!��s8в�T�d���f5k��qep9�hu{�UN t;`T6��We!��Ch� ޲
�4�fP�G(�pG_��HM�+�j�I�k�-¡)���{T�^X$����3w��[@�[s뙩zX_ɳ��)�򿈖ܱ>�,4f���K8cy4��׫|ٖ� ���������ӓ�T�l�u��\(L;��^�3�U+1ж������A����qg�ډ�����[��)��R
!B��߰�J߸���h�2F=����Kf�W�-���yJ.��{���܎���nG����zM�)�c���ۀ�!X�]U�� @�#�a(O���6;�`�*�Օܩթ4L(��x�/L�����6�H�e���#~i�Z�.�ȇ:jd��d!E.���xNȠ�4A���cW�Sǃ�u��n�لC���#+y���i�RE(^jB�b٘�Q�O��яJ=U�C��]��QVp�?T��#�s]ڗ���^����	vd�ݫ�F��}B\�B7$��b��p�*,]�&�jb��-8%ރ��g��%2�
�;bm%Xf2��<��df�nt�%	�:RP){+�=
M3 v��n6�c,?�`Ox~U���=��+P���h���~ш�o�҇�Y��9�L�����ttXk�u�挥\�]Q�og��܇�Y��r�9�Y�?��Rk0���W��1OG�*A8�].�$:��- �6Lm.Ah!��ꛤnB��RJI��8!�n�l�<�܏e�gIh���Y� ���L�o���n᨝�'�;���5&dV��$���P�����PI�㡥��a�&	��R#ޯ;i5&NS�\�A��v8Zu%��	�l����m�>j�b���/�T�<�VL���yևȲ�*'ɟ��R;|�$A��(iX5GK�q���S�*k�oٵ�+�
#S5�^s��4Rz?C�2%�i
9����έ+�8͛�o�SJ�[�9�e�_��M���/"-W�V��X��󰮄FW�}\�8�D�������;���V�V��tj��,1Z�5l�Ǚѿ����K�x�A����r��;�[9�*[���pz;�XJd�7~���M������K��ƴ)�>���+s�-<�24���=z���0��ϐ�B�m�Պ�J�g�})_#S{�Ӷ�|ƧO��[���Yt�+JZ&�;�,���*P ,(��lm�D���P���$4%�M5VV+iBܟV;�֒<�>���gd�@f�0L���o2<g)�v�����k���ٸ�|�Aˤ�{'�&Py}ǽ��d�q�0���)�bpSCv�2��^!Tùx�ḤuC�Ɓv�(����5�j#� �f�:���dH�>���#hC�$�Q,Qٛ�Rg�!�5}W!�RC���%�lͥ�+QΜ:���̞*2�WOe�3���Z܀,�3i�x$w�=����i��~`��li���
� ͅ�/��̉��*YH+m:W$�|���w��X�t������6�^�yJ�@��,����S �(���O��ƫ�Q��.�FQ[�x�O����a6!�~�l��4��s�t'�	V��E�i�v�Sv���z�d�x��x�%o��������6�S�3�](Ć0-p�:_5�ڒ�j� �q�uFD>� ��!:O�_\�����B�ju���b��zS�������/ty�K�,�`�X[�l�d�qw���ZgV��]��$�O.�B�|�?0�	^j�`3^RJ����5�w^���ɱ�C��2c!
l_�E�/J���wG�)�AJ�	��_x��܋��"մ�'n��4$���H��أ������
��&FE����<���F�.���G �z��\ӚG�x�F�5
W����e�q��-;�1l'I}��.J�@hR�p�8�H��0�{n�{/y����9�� ���F�۪W��Yu_@��.���]>��Q��:N���y��_j�-\��E�� �ˌs,�3�h�/�=��n���f,�I��0�m������6�nS�B���ێ��z�!��I4����E�LU�K
H҅��B�h�P�9�y�[0�c��lO샕s�"���hIuR��
�x����0�5�9��N�!P���
�8���M�%�Ϊ8�WS��o�
w�oULȅP�yV��>�n��R����ԟ4lS>y<'����u)2h��5X�0U�FYX�}��Z�
�R��hJ嫻�Uh��AC�3����2�	���1m�:�p{�h��M!�/��Lx�w�zӡO50���	O�~?86�jH�b.�ԧ3S��b�P�����<�=f��ԃ���P\�k*������|���1�s`ք}���3M;��B�Ic�]X�9�l�~�JO��D���|�k��u�Ĝ�Z�_޾��*��x^�u��\?I��CT�
�MH��Et9.��وN��Qˏ�%��G>�ك�������@ޕ��yPߪ��B��1�v(���hr��y��\D�/N�]�=����u=W�%D�Ё�s�)k�؅Kz��˧=�>��#���8Ӻ��?�#�������N]��	�7�'LE�FԻ[��n���i�#�����K8���E�pQ���������eܹXx
��j�jB�3�+A�vnʋC��3�](�![�Н�>O��T����դn��_�J�xۖ������UJ*���)���u�s�BaZQ��t�b�J�n��I[\b>CC_�^�Mi"z.R^>���\ �C���2��7��[U�6�ͬ_�u�t��SN?�'�+&�5O�Z��v@���j���՜m�?��<)��?jˍ�8�0t|~TB��(� ��b4=3�U�a!O{��xs�mD{;�)�{ҕ�s����{��6��mB�[��[�@s-sYj��J�X�"h�
�y��׍�!��:�.�_�$��Q�&�4�Exu���$�J{'���*8����ڪw�����;��NQ��*�`�t�!vی�〼��`�{���<ԋ/��uml�"�K�+�X�l���;tTL�j��>Iv~�M�N�<����xfSw(t����-����̤,ӝ�	�AL5k�����c�,�Y�5d���+���Y�V�mh�"|?{��iқG_�Y��3���ߓ��l��B^��1Z�[�I���,��.�TA� �ȶ��L��3&YRw��:��1��ws�I�@�5#)9�L w���$Ql.�@u�)J⒐J���ߋ���S��9p!��{@
��9_J��%X��h�U���n%29����ޝ� ��/q'N����:�a�������FڭG���L�I�x7a�?cu�<fi��Rߡ���YX�G�<��͚�'�Nk2�h�F�NB���M9	C�g&������6�
u�晭z*���ްٟ�{�c��ԎU�݃�53�(
�����Lw���>T�ͤ{�Ÿ�ew����b�&�M}��CB�
��r}��BV�߇a*�?�������c�)�=D>!���YP?w�/�=ce�>�}bn�A:]�ob�2B6�Y/���hΞ�|�H�S��r�K	�W��� ٜ�5BB��x�.���5)�E��a�uO'� n���wb��������G��ۺ��%��EA�k���NcH�/�p��;ٱKk~V��w������B6l�:�@m�9���33�6x�}������q������ ���=m ��?�d��u���ד\>�'(J�v�da�h5��[b,#)'����)U65Z�������&[]��&X��vz�^���s׸QJD ~��i��3Ԕ�.mA���}��-ðӯ�YlL5�Q�v����:��E}���6�Y]�	�V��'�F�������3��IA���P��^Ņxd����q))�������u��@�z�o�ʷTк�����!;Cݹ�ן���/M��oѝ
*j�ۘ�4�Z�֐��zN]%�$�7���������7Q[]�ϵ}�,� 2��+y���U���#���VB3�eJ�rȕ��= ���u,�A��V��<�����Q�����l[ߕ*��,fC�������d$�4�n����l�u��<����XD�~�m��U@2�̫�6~?].g?��H�B�a%|���{��״ѭ�+̒�����6�{�Ie����ZAR�H�������
�֕�;�0�\mS�+��:��lk�ҫ��f�o!���`���
ټ�K5��UѪи	 �S�[��y���x�L��������R���*���!��l��N�nc2fm��V���,TnG��v����k�_�<�I��弍 �eˑG$))�/wU篷v�^{&ۋѤ$��y&�a��IB	�}ZZ�)J�k��ݮ*[ɲ��z�����E��}������	#�Ƨw�c(�"���GVvFq�9�����;��u����[���$	�i�J2��Ol�6���G蘚�*d�(�ڔ-~�1��(���Ti���/�^�Pn����(��;^E��as�)Sj�ڪ�ٚ5|�s�*�zƺ�]�?�8
 �����	p��\�s��if#�h��J;w�ⵦ��owh�s�jd�n6A��7L�:w����Y<��fpu�ؕ�)�q�I��ot;=]�vB��^���+#��>�����{p���;1���9 �
U�Tơ"�9pOH0���+��G��[����j��bO�����4lGX���+q*n�j,>���D�V�X�� ��G�/{�����j�$0���ƿO[X3��|���zs�J���E���@���8ea�Qn!.Hbͺ�?e`Y9���#�a��I�[ھ�K�rW���U�3��J���W��Yi\�98���*�����
%��C�W�,���o�	��(����u<l|�/̥�#|���;1,C����c��!��X-�u�ծ�Ϯ�G�)��n��`S���|��&^��[�����  '�[�6fu�!����������͕��w�e/���ߍ3��̱;���n�z(���4G�?	�;�1�Q���A<4�	.W�ߥ[�4�H�zaV2u]��'�翆b�r��L��'K'6���&F�(����O$Dz:9�3����UWdƃ=��������d��>��
�KX@�ukU�q I�-wI/��){yY�����),�$�ʏ,�{��͚��uJ��-�@bA���O[ح������$�yʽ))$5q;���/�9�
+��$Cm�e�ϗ+�U�����3�$��f[�������_��ql�=�����'Ę�La��Cn������Xc޻c�򲂩4�w-7��t���4�p߈��/�u���;�y� ֓�'/)yT"ڔN,OE��j*��3Q�W�3=�E�l��E`�	����9�򇞗�;f(��ޏ���%b��ra��v6�R������6	T08� ����zW\ 0��Ž���J _�#��Q�
��&����s,}����o������&k Vh�߿�z��<S�~�f�ί~�0��e�m�*�\�Un���Y��@��QSk������B�[A*��i `�E��i"�N�H'�d����/����]�.h��
�d`��g<�s��)�$�.�$���n�jb�a%�I�!fo����U��l��_�;�Y��sI"pˌ|��8Q��D��j@�C�]��" &i�e:�{�5��U��C;f�Ĭ��hR�2�;�Zu�Ƌo�XqUG-<��&2���S��?H�+�J+O��ɇ��Ng����$>1�R�>eT���H��Td���<���(Rs78A/%�vA�q!UM���?=�h�$|���]$uGL�}w���~�bYuL� �����D��Vԃy�F�[�G��)w}T-�tT� W�L�ò�� ��Z�/�ꩨ��|
����壬tIz��)��^�e�/�<���p� 8oF��	��`��7��f�E����B��q�K�pG��I�݇qW��+i_����3��K����9�*�oZ�(p{�ۊ�W˧"�A��8��xկ{a>\�{�w���Cge�٭j�RJ��x%��CІ�'o�@������g.�Z��zRL�ڹ���"!�m�o��Mn^�phۯG(��+���!r�!z�n>?��nSw��~)������gu�I{2r�BR��>�,��vQ�]@��
��g���%����e݆8}`��֙�d'��ML�ϔ�"�Eg���y�i�.ǚ�j�r<xQ��cR=pA7��D�q)��X�3�1����[8����3�b*���Tk���Pm��������"}.]ę���%��'���k��T�>x�3W���Լ�9�좿";��x~�&޾��y����p��,F��B��[�%���J5L���V�����#�տ�h��e��;���|y*q^�9"�ם*V�l���Ʉ@k��*�o���c��&KUn��$'�e�.1�ߥ*��Ćc;�R�������TN�Q��0�����?Lݑ�l�]�*k�?pNA��.�M�	�������rN�����з:�,&*��ⷑU��������7π��y�'�;���_���{r+Q�yf廏(�ܰ�ww#��Ɩ���Z���Ú]��m@�)���ƾ8��'Q�HX�[' ��q�}��.�w��eA$�<��x��}G�p�nӮ&Q��)D�C��׌0�
�ke�B(����a־5�u����:3�t7�8�r#\�1q�=l�p�1����(�$�ƻ���n� �"ٯ��Z�ܓ$|�9�7(��d.DX��4d�
�@5N��h;K���E,�+E�p��`J���:0�� e������D�V|ƒ�Wٜ�����O������s&���I޼l����4n��d�̬�SM����G�C�\8�?�7w�mB*��a@�.�ou�v��<_F1K!�]_/g	������[��ퟰ"	6�qi������[�|�푹3�N��B�k�3�iu�r�&���R� rpldC
�^F��,�F�H6���b��2���]�V��Ǡh�\�!V	�����L�@�,�I�sE�{��C�5n)����;��Y�~�&+��<�y�P�܃�E�-tbCq����93���F���n�L����_���y��O?�(�	�ͯD�8�/_E�3��8ZQ��`�d��x�mI�L5��
뷾Qǝ!.����K�ѕYS��2�������Bo����=��a�2�-�)Ub��I���.�$26I�����dŪ��9L%�(��h��_4qG�>�Le��$�Z�;�����Q�05'�ᲀ�[G\z�dfX�\�T_���%#�)������H���q�.�v�8�~
��x�о�)$b��:G㣐�|���.��_���z�e��ZB%f$Z\�|S��g�L&��� m�ߔ8%����E�J����<�<X�H���8���:g$j�T�j���j� `�s1 �9�[�	)q��@!���;9�����+wT�v��"���>e��(4�@(�zL�r�*��U҄�F�FTn�>YՐ����Q��TeC���Q��`F��8�$�yK���ؗ����	�PU㑓2���_+�#�[e?�7*C�Vid���fF"����!����c�k�+*����\���z��X����ɦ�^�8mx��ʳ�]D��c.�vG?����ۨ�xnnîg(X��K1�,��0.a��m���օô�;>>���Nd�K|_,�z��6�gA�A6�8i�ŝ�وO	l�U�&"Y$niݗ`�3Q�L���9������ �r0b�ׄ򧿄2�՚�YҦ�?�2\)1ɕ͜���8$�M��J���y����ԑaާKr:D[����;_���-��Ah�E�����g< "mA%B�����ծ��N/��}����ʢ"U�-�@Յ����m�(8w�S%�TT�Gxy�D�Ԟ��I"�|,	V�8�I�!�8��%ҿ�m-q2��0��@̝��������W�{[A�2�!�-�,'r��t[^��[���(��k�	����ܮ���E^�Pa���
��Ϥ�Ptkԥ	Ի�E�%(;[�V~�	=�x8�R��b�Y��1����Ǎ;eZ
��̩3��hn�"c�Q�k|*�"�7���%*ר3��uf�*���
ε�ے�{�����k�=H9�D�at9c���_�PKl���9i[�f�)��ۦQJ:�4\�p[�c�K�A��!��˥5i�g�:�XFS�5I�;f��eh7"uy�ïЋ׈R�h�̘n�m�2�Nݻn�,�����~�?�T��9Pni9+� �tX]&��v���^�D��d�t�.7D6:�I��v�pJZF��L�HkznV�1�<(S��=�)�S���R�+��ŧ�Co���KW�\�a� ��0�⯷;����g�������_�Fg�7�GU�P�N �|B�M��z��ˢt���Y5v�9#��6�0>������;�]%$��6=���QQ�o;>���	!)n$����X/#S��y�_RV�6>��r�;���y���8?�����t5B�#���G���j�g��^A�_F�Ť29Qi�}�r����6��g�%Bu�Eb}�ܰ��Q[y�k"��Xʔ�����7zPu�"��&Dxy~4�E[����;�X�e�̞����ި.�I�E��"Bʕ�����¸�S>��R�>�ir �h�۝��U�]�"c�b��8��t�ՙ8�4k��r�z�!�Q �*ڀ	�$�p�q9�/@BL���:�Ԏ���NJ����Q�pK��Jy�fTVaL�Z�%ZG�▊I׾2�_L�/�*n@��}�)��ID�Ȏp4L��%�L<9$)P��ܕ$J	�6�[ì���o/�y�+���`�D������%�����\j��,�����������N���!5���X��������0�4��u���R���I�g��}Z�W�mᜁ[VF�3�pGS��3���M�Xɵ�?��W��	D����d���|�p�v*'d�w[��x����M\����l�ѣ�?]��mg F�h	�����^�b�'�1����#�_�e��XW��9~���YLQf�Z:�jS�rC=��آ�BG@YA{~��-'<3(��(��p1�e5����۹��
ǀ���6y�� ��?����gq%;��� l�	��}���7�BߢV�ޞ��#��׷�ω�X����c�3�#
 	)��㆏/��~��$��#N����]D�K'����ȟ'�&�@�$?���8߾uE�u��/��d����G�f<>�-�%IH6��t���KZ��u|/(�(s�8W���y����,�����aU��sv������"
r�*�ڼs�iR}�9[L̫=�l�\��^ko�\���>��(]���&�O�6.k�qO��6}\�S�{��5;�y�U�-@�>�_�'�� 6D]z���\�UB=|^i��E���zY�)�y^�x��
����o�k� ��L;p���e��5���;�њn����h��i[/r{͸6u3.�D��đ��#Ω���1a ���rU�+��B�IsA֗��4>`X2?^U���GM�)��T�A!�1bTV5c�ˢ��e��z��X����N��:J�@{����GCOؖKS����L��X�[�vL�v�]��.}C昛ߧL�RaTE�I s�1&e�ń켐4���Z��߳|�������&�-�H��9k�%�{�@��λw>��҉e4Ĉ��� �o���~X)6.c��[E�����6�A�;f@mjC���DxN5�<-#�)�d{5m�������g�Z�������I�V�e���0�.��[L�:�G���VO�Q�hT]���7$�GY
��K���w��b�~3c3�ξ,�
-���s���\��3h�� R M�����|���*J��rl&�jJ�?�)4$�Q��+ڥ�,nf�"�'��!|,U�h��I�N���2�������a�1���{���f��#\�^*��e�m�g2����pz��7�Z!Z#܄w�e�IV��(e���������t���1��Y��\p"N`壜�H������������,��q�|���,�)�u���s
�rw�ѵzT����N6��B񴦝Α�Ď�X
���L��K�8$k�����X �۱.pv�R�yZ�� +y bσ�����s���<O�\��=Y�+�Z��eR���ٻ�"��8�9��qD =]��5�J��3M���w~6�Ne(G~��9�����N�NIV2� �໺m<�zօ��6dHN=�ꅡ@�|	�4{�F]�D7�����e6�ޟ)��x�tֹ���VA���q9��-��;j|d�p�����ϟs�jP��j\���W��2f�B���2�WƨÃ�l�w�.�üj����v�i��+ˀ��͓ɵ}��Z�	
Z� >�	���d4tǢQ�'Y�%29]�(�#�]�׎xLA�ć0�ġD߱c�vyK���b�R��)��	qQB�hg_�|�=��yR���ƙx�ߌj1�YZX��;�ݸ��ؿI�t�)��eR�s �O'��V석�@���<;԰&s��~+;r��{�D�Mpre�M󂛒Y��A�M��1�{/"k���A��Db�W�p��=��
}��F�ȭ�����G��h���oW%�Z���z���}Ώ<Sx�k���	�\�&���3���B���p?%�\S%�o��Uy��������|4�i w=��A,�U�)���<Vo��8jA"m|�������e+������K它�mr����Sϯ��VS9\���^�^p".���ς3ߑ��0����<km�-8m'̚�o���E6��38dq�3y��յ�B{e�@#e��G����_���W>1`���m��R���w�C��*�t7K�	�ฺ�}5� �ԿV���t�!��re�|�aZ}}Q'�_����!<)�ʣ�)X7�����1��`�����dִ��������� }���M��B^��Y������Γ"n�v�d}hk8��8�s��� ]@���3�������~�fw���B�=�;[[����]��4Z8責�X�U��K��J��⛞�'j�<�+��M&���!�
�^�IO���X=\��v�i@+�պ�`m�h��?��(�����r�`�0B�,�粸11^��̩Ș�T�j��Ď�����Bw��ROt����x:_a��ϳ�P�Pcw~U���O>3���珄�h���VO �2�NK���B�P]3cWԨ�U-���U�e_b�\���_�!���;k����2ױCN�gs_\�*O̔����o���&�7H0��0 6k����!@�k�I0c�!��"�o�$c)���R%; �D�}�3>�C�[�IԨ������5C��D1F�Vc$e��G��_���/Ӽ$�/H�r�3�<�ίަ\֜�ֆ?����W,p����=S	C*�P�c����X���N�r�b�,��"�ktꡫ͇G0S��<>k��pL���yD���Ln��ӽV�����2)�Ev^ө�CVE��'���G���촙#�,n���扼�ϑ�Y�+h�{̮UȣEd �U��
y ��?�o'���8�0ee��'�Pda�x��H�Y�G�6�Ӿ��č\R�VÍKr\�U����2XW��w��Vcɍ�՟g�WT�8ί�T9q�¬�X���N��ڧ|v�j4���L�;���6�}�U@�OԨ��Dky�A�0��N�d|KX���ů�i�ֺ�`�mj�+p���O#��x_z���0L}W����I/U���7�79�ms����p��W]���~�sb�,x?p��u��i�M���������
�2��Aѡ��bP��7�I�=nl��'��3"�E��E�Ș����J��gkpUj�X��b�2�x>^�)�_b�E������8��{B�qZ��~v��� ҨD�X��NE�K��������S��׬��u��}{�d��󂦞����@�l�K��Z�����>��?�.?r��H��$��o��.�|�`q�j���X<pբ���qǍь9���U�Mw�(UOAlP�ER��+ol�
�����iiZ�MX"Ԧ�e�F帯�pQD�q�G짒��=���,Qӛ�d�8,��=�?��~������8|�vhݖ٥��ł&�����.�A��!�qK�F_&�B}�c��%��D�'R�3�;|���uu��p̺3��v������Ox��%�s�ҳ�/�J��w�_\���ek�e�#Bݪ��o�#_l�16�F���X9�ݮ�:v�6#�?�_�� ���Jݖ��K�����rr�ª��-r���N]�e@��Ւ�LexR����I���. ?���$]�E5�^����;(k�U`m��i�8n1��V�L�9A����J8M�#�H��������ʊ��+g5)dgp�qe׿����1��j�Q���8��=.�,u? �cPK����r���#��� ~�S�r��G�(��� !P������g�=�r�d�1�,!o�Co�/|��'���3�@L~@y�B:��&�fr��d��	��v9��Yx@j�����`����9��*�y)G�֜lg��̧N�2�6�T����{^�Q�w(~.��[�i�V����1������B�Tʨ�U#�D5�~������g�Y��>�bz�R�!�6U?K;d��~�5�#I�bf�~ژ����b3�j��o�E[$3�
�^���q���v6㥌+�m�N�ٔ�u".�k�/J�H�zO��wh
��H�
N�?�^��.��	�ܥ�k6fΪ���Q��7^�a��6��BS�4�����?�p�y@Cp� �� A�sf4�.��O(ם�� �D�����7<i�̏s���E[��Q@3�N�����T�?�x�Z{���[��3���Œ+1��{��ij�B\8c�L
�.�%�2��j�V��[߽�~Dx�P��)xF*������i �}~��=21~�=�˹+��5"ѭ������;��"����>��y'�DZ��A�D�M�q�1Be` n�/W���R�5�J�М�X!���T�Ra�4Ѻx��ꓥŬ�,�����F�/�E�!��w��[�u��a�x<�N���a3�Q�AE����{�t����w#��w����ko�G�.��� ����������!xX�-��ͽ�����;g��9�3�U�UO=5�{�wz9ƀ5'�
�+�zR�`{Y�v�<�4��7�*^O�&# E����j"�}NSQf�Th|I��1q!�z��}X�j��%���H�u_89yP>��ф��Z'��n;���
"���ï�c��D�xx?F�~����p߬�����ګ0�ɕ5|�cڎ/������G��^�H��Gߡ��YR��qc�F�)�a@�@=c1�8E���A.I5�����J	DD>�Τ�^��ly��xJ�;)���n��h�=�D�6J�s��@�lW���'&eeT��+T��#{��	��a�V�M��.�Մ�����j�~���-b}��GH�0�xv󙽦��I��h����O�t[x�&���9��,�%��x�®�"�~���{��H��o#�ѣ�,4�z�"]k�D%e!�7�_��^
5��)��SOR���J�C��p�7j�.~��Aɠι���8V���_Á^]u�������b��<v�3I���9�#���\w1n�0��vj��t��~
���u��c�tj%��TH7��c4E�/�M@�&���E��a�V5{�9ts���3H�քb��I
`�Ĥ�7k��*�5НV�)+(��k�*ѱ��t�ҽ���֛�w�׏K�RTt�u �y1S�\*��v6�@���&դ�c�~�漕�/��*c��v9*%�*�p̋�mQh|��	���3~�Z���`��Q�⒗��G�W�����D� �cHh0����0�^�;���I�y6�C5�dL�����Y�����I����y��7�}[Тj|<޶��;M5�a��~�Ѓ"���o���.+ "~��&�ξ����NF3v��]R��0�n�H.��Nl�}�����{q�Y�%�ycJձF	$L�v��]}�ԥ�����,�-[D4V��	�j��E����ku�\��n��hf[ڞ���:������]��<�\�)<n��B2}�d�#�2��/�$eH�u��ȡ�����r&8��ʖd��������Q�Q@_�f"�".�Z��$(!���2�H�N�ܣ��|}b���s����K^��
J�t��Ũ��,B���pXo1� ��SNѵU���{��]洝��hV ��~������k��c�r=F������.z��,az�|��'�k�Z���'l���
���	�Eq�:j�	�.�l����-=����� F�����>���fF�w�2�d��M��[� =��Z� ����V�K/e��IPd-���z�좕�N�\ű*ш&�̘N�ܓ���o��"I��N�'��NKe�Y���FkWb��F�������ܷz��9�����߇}�(P+2�9��4:pe�a�|r�]���;b=�X)���&�;T\
���E	R�;qt�	"�K��B?/ ��!���-9|s�\���'dK^�vآ�Y9�A��2͵�dtFN%H��^̝�|�����.�IhT=��/"+�F��r���x}h����2sZo���N�ϦfO��EU]ŴuĸŽ��1p��HZ����.�R�9�=�giA�jC��~!Ti�Gf;���fw�Ǽ�Á�	ϐB�!��'�:r��gH�L���G�X!3 �ct�s�2�Έ��k��~7I�8��-
��De��t��k�S�}�&I ��ɩ�V8��d�ЁI�s�Υ1�x�\ J�Ó�Mŋ�*"�hc㢟�	t i|+��"-&�;b�v#�d�x�`�*�\���5umw���_��WŊc8�H�h.f���>��ަ�ҝ�Dn�c ~."�������L@����%t��V����Y��i�3mtϼL2�&7`y�%NlS�����S�ei���j&��-1��i5!kTZ��Kz���[�"��^Yף�]�S�M�^��E��#�Ǌ>X��<	��Ϫ=�!�6��"�!�n@��m��,�6ROW�&�8�'����3l�yˊI�}]�2A!��+�[�e�54��[%�q������-�+��[�lg�5��(ew'�Ѱ`�qF,��l�l&���[�L�Q�����d�귗 ���IӉP�'�TX8�&ކȥ=�p��"�X� ʬnUE	�cl��m��B�L�l�(� ���wP��}e	�9WJu�֟��?�~{q�C��Y5��V�H��$f�?�gD����3��Mߥ6��&�Յ͎�܏m��b5��y"���h�8A��;���������u��x����-�i��WI�I�"*�3�P�(`-��g"�;��@3���\�=X�>���cB�U��X�3��N�9Nb�,��(�/��z� [ط7=���I�U�vrq1h.㸵��(����w0�d�]�/1I�;]wW������Jp��1A;&�زN谳����j�"�V~I+V���X�2��������X�ҙ @�s/2c�����6zh�&Q��(JƐw���7x��F��Z��]{I���sfxQ��)�s�G1zY	�ʉ˼���戔L�G�Z.cJ�[=+	u-N��L�A��ߞm�/ݝ����VZgJ*4���)�b��]�j�
me?tU��!B��C�B*&�O���H�x�� ����*��=ƀUӽy�<�w"5��&Q�a-r�`�I�vr����ɖœ�z��:�л)���!�w{�\AD�yq��/��
�U��^!9n�=wv���{�~���'�cMb���"j����(	},Tta�S�SĒ@��&#*F+J����e+~h�?�Z5\q95��¯�ە��:�q~]��O�~a��3�0����\��	2$x���+�R�U��X��V"*���u]>�
{�������3ZEr�@���kj�@��f�{c/���Q��K*�l��$Yʎ�����t�2�	��d�ȗ��͐w��:��z�	���ڿ0���s]�ڂ#������#�C%O6.�n؜���j닔c��o��;�+:mR�E�� ���8n����۶O���}G��#��Q!��ؽ�Q�����u�y��<��X@��T$cy륜�	�	����يz�����'u(Sڼ��a!�?FX[o�Li��h�X�9�%
���s�H����m=ӣ��6 qY�2��`ٷ����������h\��]
%&�J{�d��0ӯ���Z��~I*=-��!%� �y�qS$
�v�ƎP�ܲ�<�e~E:�~�P$(�٠�C(�R��g��d'���[��}*��ې%o:Q_z���|NH�����	����f�9�o7�M�����l�#�<J����5��֞1Ѩk��6�L��i7Ǽ�f�Dd���z�p�{cƅWQ�z6Y�t��?<)���2��^p��ڈ�*�N9N�M�C-�n��E��z�r��6�)!5�TYc�GՌ��B��x��ӗU���F��ĥ/�n[o��tD�#'#:�2�5�>8!*�O{}��ѭB�j������P�ɨl<yڜ k�L��N�TV�,�Niz^��x�_S .��n��7�q�V�V�>��,E�+��y�f�nZ?".d	P��^/�RH@�l� '��;�ʢ*Ey��}�-����Š���3Y�����n t6̐����Ҭj�IQ~e{X�^�g����k���
�tԧ���X*������;��wK;��A~�Jĥ!�k���xnA�@�5���iIǭM�1��Õlj9�[UR��z�s~�G{V&��O�d.�T�b�i�RE������߃�\�A�]Kx��SJ�wE:�l�W����[�X���Jd�'mmI�Z����; ���ZQbc\��I?���죑Ѧ���j�I����Ҳ4~��~�{$���<�_&�T�kw*<<��t�R�^���.n����<#< �?������\.�t����<o8�߻�l��Δ1OE�XN��R�9m�� qusl�蘭/V�;��a����S��z��*�Ё�l°�J�Q�aw�٦�?�y�u,�IԱ��6!C�_�s���M���}���No,������J7I&�}����)���������O�ך�z{{���uR����!J�[�Ҝy��z^�+|x�F9�^���yX�H�T�)$�s�S}"��b&p��)N��[��O[5��U�����A�!!q�7Β�$Yܐ��ntr�6�/~KNP��f�N�r��_at%BB84�ar-�h�s\h+	��� ���x�b� ULm�����5}o&�}�0���V���iQd����**��x�ՖD�D�)9�k�*���'���/\�a�DB��)D��a4ro@Cvd�)�=���k)� �LeL��)2�rȌtO෯	S�����^q���gb"/���0�����PV�w�I P��sӹ�͝�{b��*A���iWSj��c��������?���Q��9ƺ�;C��|E\R�?G�W��_?���`ö�P�J#�=�#V�x�n�Z0��A�B���e-|7�/�bz��s:�n�~1���gZ!��e��z����|�2絧����ԡ@���Ũ��*��⢤F���Ϯ-���)w�Y�d�pm��J�Y%�b�Y�����4_�d̸!�t�kf�.ۣ-������j����ķ� �X<X��W#��== ����%X@�d?t	]�"Ԓ�IcGȝ,M��A,�m#�Rfʅev��sPPl�PE�T�I�C��O�B%V��s���ӱ�/z��:����kX��kQ����c���ɹ����$������׭��{<h���G���yi�� 1I��~�F���䄔<UtK���?Z��r��fu����Т�_�S'�g��B����:*/o�l�r�0B��9"P�Q�N{)���?�l0�u��"�j~w����Xnnnbq��@��uA��"耞!�o�XN`�+0N�^\�hӄ2�`����)f����m_�S�I|8�椆�xԖ��@C�'8Xأńu��@�^Y��%|+��g[���3M�NU�jئ�t:{]�2i&�\Y�4�xK�ēf��I�@R��t
���ER��o0���|�e )� �C0�P|��G������$$<$o�Q�Ż�E��1ƅ��J�ot���T-���G�:�m[0��`��~I���vw;�ë�`K��W�6�$� ���q�tNӢ���ǉ*O��DS��2H+��q�Њs�a
p����-rQG}2)Џ��{ҷ�~���oΕ�t�Ǜs���:�\�qt(�_�~8�~�7�ě������c���G#� ��	H� ���K#������2�d�Uu�����B�/�?�ʣʫ��p߇\bY�9>�a�LF1�n�BhbSڄ>E�RQs3��Wt!ER�$�D����p�ˍ�$s����n̙�\�G�$��͠�#�Grɽ�P�!ִ�J��ѝFN��@�p�0�Ͽ*CϽ։�g�ނ���v��<��gP��	xs{����fo��Hl�A qsޑ9fٙ�仙
��׏�
��:�	���7����$t�~��KF>7�?����H�Zmre�_�0n���T�r�P!��XS�Tu|�ݵ2ͩ���P�><9��Ka$vb�!̯��.Jjj#���Z�A��D[�X�����j=���ƀ+�-�����U��
���Wdܨ}�6�5Bbb	�{9T4�8Kr����۹<5J���^�q�2�<�LЎ��Oc2-{��0�p)��'O\�(l(�i�N)7��Fyd��ۯ��OCeP'm�����[�	�dD�t�:
#: 2����/�p(�*�&^����x����� �R������IX���.Ѹ!���v2����I�/�!ſ��&�+u2�ϳ7]#PB��6߲�Tt-T�K{U?,to�L��P�����;׎�R��Ԡ\�r"�Pn�<��%�"���R���d& fRɫ�#�\��2��Nk��BGd�:�)8!���+IY.r�c�Ǿ��L���S����/e�*hI�H�U��b� B&;(ӳs��M�7���,�V�V�����b�h:!>���2���Ԋ�-���LpD��S�H
�r�H���V'<Sp\<ɣ�-� 9H��³dUck���
�W�M�p����<���9c�a�d0w!_�B�_)aB˖$��o^�(��E+ۙ<��I��IH����YwV~�K�@@5�	r�1gH!:�%�d���ʀ�^�L/�h)�
�� U��5UMj;N���e���Mo�}��Ao��]x���~
��	,���o�Hv4xy\ԡ�I79_B]8e4��`��D�G����,v,�B��������s+йu�[a6'|?�I&�����l���8=��5�܇s6��	�y^�b�U��Z4���
t���yytleb�-�
 ��=��̅�T���x���M8�~>�;.P�w��9u�]��ӵ4��7K���y[`Vx�f��Z//��Y?�E�N$j��m�y�!�!�FUMF��ݩ�KX����lĭ�00�7,��^()�<9�L���bJ͗6nbee�>���HŜ+F�tCl�q��rţ�KrV�X�ۙ�7O�Ã�]���^2(���LR��.'�����!N7&�Z��0��s+~f!��ވLi��M&'�����a\S�5�3++5]w�P@�@�T��z��&u�(_r�H�q��~w�u����sZ'C$r|mb���J�T�#��4r�<C�b����IQaIQ%f��rf"K�%���l�ħ�j+)�)aե�
gp��YB����dr$r2~�.���Z���� "��;�6����@��o<�u�61�~b��q8�s\����w]����G���@2�%�(��}��V;>G���;��m=Vc��{�?��J��W��ZPo�d\����,��m=i�d:(x
8uڱ��0�H����gʤ��耥�?�j����g��w�p����������<#\6�����{�Utr��V��J(��#H��l���^���N����4\ΫWd�p������26�MZ�b�oK䋭������9j��kf4��'�Ϛ�\ٟ�Ƨ]�ܓ���l��t�ʚʥ`��~y��K f�����Ï����W���>h4 �7ig���wz�>R���e�
a�K� ���;:ɲБ-��sN�-�Q��!)Tp8r2雜�Y���5yHk��f�{P���&6�-J���׶��
J����']T��!bO�!�()��o�epo[DH��頂���a����>��১�����<���<�e�j|��J���^hΐsw�jV�P_H���&�H� �=z �v���2�Đ5�R���/�^8�G9��>?�K'�``��.�n??�M��w��I��5�&o�*,�����.�����`I��@����/g���m��',T'�`��=��D@��#���+�L��hI����yޞKD�s~���'�x���@y�Cz@u����^-,�L+Ĵ�rm{s����;Ԅ�"��,�t�7���ű�|@^�v���5�t�Ci6������Ӂ�%Nv�	0�H�4z�e٫ /����8��"�E?�P¹�Aa����u+�L;�_�*��DI��D���W1�])2쭒�ESn���ěs�W7 �!�B5��M�H�2-��<ɦ�G"A�GH�����"T0��r4��ċe{Ъ�g�����/�e|�\Bԙ�-FUx��Z�A����tmĊ�G���/0C`Ǡ�7W��T�Zk�+�N}o�?�Z�0NIz���":_��D�<:}�Z�	��+:W>��_���+7`�}�ъt�"0�m���Ր�
n��^�{q�s��)�u����(�?s��^v�Q�W�w:���t��Np��"W�Pe�Ė�JU�p�nx<q�����ʛ�(�Ʃ���b�!qn�ǃVK�OJ:�� �8����bA2C4i��҉E��k�Կ}�J:m]����W|���;%��i���bN�5y���L9�/���qd�r��8P]�>�r��67P�V'�;|%rMv�)r��!-��"�!`Zj	k�r��1y��s}�b\�g��S�p��2
�>E�n�� Y]�p����I1y�A��8���]���⾻�~�����_��>���o�n���_z��.�5K@3i�+���iJn�bs�5����.��ʙ�	�)v��!��<���>�e��[�|f	I>��z�)��Bl/>���Y�GW����w����̓��%A��ia�H���8����kT�6t6}��sА7�,*6	���e2��$� e�����WL��c/���fgj�da���ͼrA�:=߾ȫ��/�|�L����G�����YB��2���5��
I0>6�f��MK $mӠ	��Hi�F�*&u���6��ʄ�Df3h0uV�CYJ&�!�9��i����2�m��a�'�\a���?�SSk$0�h,���hv�[u�3�P0s�˅3q[���d��k������x�2N���hLZ:*Ps�!δ�Q�9�Fm�/U!�^\�.n,9���	�kR�EԣW��vy�a����>~��Dn�]��'�n�x�``��޷����P?�=�In��kH@;�Itm�P����dT�_���O�<?܏� �Ǝ ��tن��>�����t�>�|���On�}����](��]�^�!���Ho���Y�Y�>��|�6ْroixO��4΋}��I���:"Qk�
�ti%�c�4�d�e]<�k���>Wc���$5ݐ7�B���?�R��K�WR%�8)#ƕG�/;�#W�[��/'
�hSWE0\*f�Fkl����jM�fr�c��8d7ʇȚ�RkH�]»N��!�����7#Q�aϑ����r����ՋV2��!��5�vq�޻���pOU`���h���������	}�$W��L��W��	�2���lO׬�ɞ�g�E�7F ��"W-,�f�/D\�������FyrE���Yl8.�>|ivݮ�	�������`��C�3,|������}��:���|(b<%�.��&"�0��_�.I&O�o�ު%W��­B���˕��Q8��z��A2���j��PP���(e����WDo��!�Aa���л�� �qi۶)/���	&<�QJg��Gu���UK���@��"�]�Ԏ��L����*T]�:�+!s�M�Z��O�����t�o�+7Z}w�yhp_̖�]7\�p��d�Nz����6Z�X��7��f��zN�Oǒ�DP�X�r�>+����c2����榧�ű��G���v�q��S���~<�ag��f&��
��V39ߣ1�Y�	�o.���N���r�;~� )밑��D��o.�:���g)5�֩f~�i��
���|�Y����uEB�|>%�Ҳ%����(�2<���	E��q�L�������q�S�v�ͱ�;��Q�rR���㢛=JR.�T�/�:�������!��c�>�ڗq�>a!�C����D"ޔ�ڌ��xJ�`�?B)�9�=��^
�]yɎX�u���Q��h�y��~'�7�����8oϠ_�I�jT^���{�o1���Ip4�����Ӑ��$>��u�[^wH�
;z/1RvL���"O�ЫC�0�L�r�'�r\w��8�<{$ĵ� :�|�}9��y؋�c]b�~5����_�G�Y�U�^�t^�"e�h��C�Z�������do��ŨW:;OT� ���G2�(��koJ�E�
��D��nw"��dP� F�P�j�?������pbF�g��a'���$����@H6%ca��⡅!r���M���߇�a��7�j�Ce7�;�!*�Ur�`�(�T�, ���ыjyvȈCxp����� ��������;�	X�K�<r�o�����7���n�ӓE������ˎ���`Zl>Ro)��[�',Uk��&�b�ܝ_��b�a�n�Gz��4�~-���W�Y�%Y�y���C:��c��}����x;������2Iw���E:�}��
������AWLC�,��C�����wU ^�*7.?,�%�/����9-��Ӛ=��vD4�;���ᘒ19���*N�C	�^m��Qé��vO�!�!S¶=G\��D\��M�f$o�^x-�{�|�L�l	������R����pщ�/8�Z�W��1k��/��qu�b�r#�9�&��SC�E�/�W�� �垤\�λ�s�f��1=���P^[6#rZH �J���?&T��lO�:H�&�,�cY�3��j=�"w��k̌�*h�=�4��>��Ӻ�I�G������Њ�f{J���eP�M��p�3^^�U�+:�Z��x8��l����9e���Y��� ͓g��W&�����4���+����-<�d���e)[P���'�+���)s��)����X _O�ayA���#��O���H�q�l�`f��u�q��L�����@�j�U�^y�-/q���J+k�<N��h����M��4l��B.0�%��bUz�~>'�=�]=��h7J)�za���N�A��
�t��U
;;��T5A� �=��$i��.��B�[K��2�&�u�s�P=2~z�<$;N��m��B�ݎ���	H��!76�w1$���?"�]�?�[�/a���.V6�y���� �;������ �4���D�M�p���_qe>��~P#Q��CE\`?Д�w��#����Mv��N��gc��Ƀo�i뵚bZ�_p�y&[�(�#5�:��}u��	�S�c3G��iW%M�7�H_���D.9]�;|~���M$ ��7���h���{"�}q���e�-�5��*�����$&�9+>ynq�2�BM-��mP�1����{��?�=�,�0���lXwl�T��������iҡ��<����z������V�p�j�#�=���<�MaޜA� ����az�i�i���i�3,�<�~q5�}�AZ��l���b��-iz�N���\�����G����sXÓ�S�Z����1�?iI�����}��}����j�*����L�ڊ���'E�/�-�P�"xY'��]���W��u.g�b��|R�ݨ����|��Cͦ�q��8�z�TL��_��"qt�pٖ4���^e��x��G1��(7S�R�{��{�jgv%��"�c=�b����SBʵ��b�:5�6�	�?��V��+L2{�=�X\�9��9�o���a�pr��+�~{���^����߰�1��Ѯθ�}�@�����N]��I�>�p��T?�_<��������fe�lU4����Y(6�a��5��/1u�\�1�~%�a��&}TmT�pڗ�Ğ�-8�:���1��'t�K� \P�'��3Ol>Ѥ�Q۳����r0��3��0V��������	�	��,�yqF�ɣ'��యm�.�����R�^Sk�3d2�GZ�
��`�#[��}�=�\�H ���,/�dD��ň�-�:5��:Uc�l���ǧy�2òi�����O1��[�X@i���̲��q2 �=���E��|�'�<1(���l����Rmy��'�^z��^�6�����:�r1��2��.�BN���p1��.>R}|�ک�9>n3�t3�K�]8��E�@��QB^��Dxpu�À<��8Y{3_��ft����cp.	o�C�'׃Ԕ�Ka���Z&�OԒUPR���&#�t�V��� T6Bg�VT1����-pmh�u�+��	p�"�A�3O�'���q���&_K�5\z�����B�cZ�6��eSLr?P�Q��4�6j����DƆ,�Y��}�#���������y�ޚ�:�̄�?�6���.�o���yt����ɲH8��|ln����W� �^�ij����� '~��x�7��*tqN�JfN _f��Ӭ(�	,�>��1����=�B�C�յ�<�tkH��p!C���.]ш<��?��$r���"F�a�$rS�d4��n��w����Sj1�������+�}��;Ш{�o��
�0U���s��x+RZ�XY,��5��i�T�xU�Pb�)�\�h�cTmj��6	m�i�8�|��c@~uD�J/�p�@�&�	����.���"� ԛlG��n��{N�" �`ʢޯ�"����#}_�H��&?wGU�>z��B�������SR��&XNr��ZR��p1}���~�)��&Г��G�C�)uJ�v�tI;�)�y�TP!�
*�¿?D3N"����v8�nۆ#�|��YEGG�yoT3������@�I�/���ˎn9w�_yF�:I ˁHF�ɲERc����I��8 ?���EV目�@�La���S��,(���v��J�!~��$���/
�;�K�l��l�N�@ٵ�(`�	Қ7���-֢t��]#6�oW�ψ��SN����g!�d[������,MD�8oCd��B	��x_�	��0���bU��'����=�Qߝ����Έ��2��)N''K��{n]��A6]�h��lqLXU.�?��P�>�zm�m6C��;�˓"q?�)]Tp�xP�p�.�@C�bF�>5�-��*<���x�� !$������I�������)m_�;���X��:>��~tnG���A������~=�1�ZL�p.{���S Lj܉�������J�e�S�*��a����D�Ad96�F8O������/֙�eN��w�$
�O��»#�[zK?�r�� B\���p��������nvx���>�"�ދ��c��'1���"9˖6yc������n���x���|4�,��g��UʯZ!W:GU�ںެf$�J@j9W˨���)�v�"=%��Ԗ3zL�x�;l��0wO�H�L[�S(�7�*���{N�i��+CD�ۊ���ㆃ����؞�Ż|x��������;,DDN�<�� *�	��BP�1S T4���e-E�-[b#?�1�6��(�#WR����^4���b@�C��Fm�d�[<�ĥթC-UKdH�KJ���'��Ճ,3l��!��co���C|��AW�*���1��뛒6��)R0�)�\�XK4�!j�<�$V$cQ��e;�;�-P��M�Y6	��	M��F�7O���
W���5�[�����k!�tB��������c�;��!��r�v�����V(F�>����uI*i�=1ک��>:g�g�?�ݟ�y����Ʉ�PD>�@,>�p�8��܇#�9��3e�a>r��.&�NP	ktw�#����%�\x)�ՙ]_���HA�O�}�!�@��Jk����8[�/��Kez�g��v��*Tx����9w��/�}����-ꇹ�,����:�FE�!�z�w�y�)�@�x:n ���܎���/������M^��oãG�����?g�����9���[o���#v�:aZ. d"�!�$:Z4ᓤ���(��N�ɠb���sPƐ`�4��_����+�z\<��~�y�9˖�wYvf�:������$��4K���p¥�!K{��T�!��+{#CL?�ps!
��<��o�]א���s)Q��c"��on��Ҙ��L����!A�!�?P�\�m�C�)J�#���2c�y=����C޾��
49�O�P��]S&�#.��
���*�>xM�O@�/)���u�\Xj�e�u~��.��l��\�!`�����>)N�|Z�ac5��=$e�gG����|o��7Rt������PX�-xp���xÚ���Ư��I���\��+`�bB��*V@��F����FS�����.��K���z��Q����',7���MC0� ���������'n6���×h7����j��� �'_>����"�L�N������(����Qf7ï�ߊ"Fu���sL�4��H�ơBfd?�.4<�N��M������D� )+'�Fp��N�� ���`4;f+;�L���l��C�݇{y-E|Ι�p�?�L�B����O$�s�ř�_�ۘF`�]�.�� *^(��c��hf��C�Bd� ���05 H����CC��6)<1��� x�}��U����_[$S ���R���!QzJ�U���Z��v��9�S|=9 ���F��it�Y|`����{�+�E�J�B2�i��	{!�
uVL[��W-��f���X�43U��0:�@m�S�m<�2[aE�?W!U�r�u�۩��"�?��,� ��Z��S�xl�Dm���@C���1S��طM���t�0�l��Z�R��Ц������uf��IU�~V��\J4?�����&U���fr�����2�9�.�[�k���B2�#�+�Y���E��rx (�޸�m��3��4
�i��q6�0a�6�\����[�B��*�P�����:)��[�!i>�ã��/����B�_��Xlf��b�Ji���`�<_,H� U��-6�&%�9��y��P�x�S�
�f�}�TRLcl,k�*�n����~8��H�_g$���x�� ';�Z'{��2<�H�;-2*���h�-����=v_p)���c`�u`<����m��p�K��@~���4A�����^J��4�U�~v�`Q��PxWbR�mK=�� ��9oRA,îJ(�,ܱ���W����FF�c��@K֨����ql�!o}�2)�Ps(��?�uqv���^���3���؈���@��wN����@+e�Zlvܳ!�
BIͧފz����}i��� �I��
 ��� ��}��$ι�Ko���	�J��[��W>1	I�����~ǩA�3U��z2KvE��F+�2Y�aǙ��	��f�u���y/��O�YKZ�����f�d��'��p�]�N�s3���v�ԞYՋ����N�vw��n	��n��=��u]�5>�i\��V^V����LŊ��WH$��ٝ�O�<��k�7�Ӗ��D��d0Е���.���o,���!�8���q��^u���x}�ﵿ����Ns����:�&�G��q�1e8(�6Q����^Q��[��i�>�I����'�ȑ܆s�QO���m�	�i1�mz$q�"��|�h=F��j��M<ᛯ�<(��rt �32$��Rx�WfQ��n���_�[:�Z�Hܕ��?�QW��\uz��-{������"�n��k(�߽�_p�|��O!��� �͐���3G��ei'^���S����l~�lEL���t��b�}�xna�lH��}�r�����d������\8�A�7,�`�j+����WRO�M�P�.d���Ɲ^3b�-Ư�ך�ڧ�zVr��$���ﶃ[��#^m��BN�;/�x��Z��a�x�:;�t�^4A/����1hD&��Y��ux����x��.�^\�N%yG�s�"J0�C���b��p��!������[\�#��j�r��e�=edB��;�	�T�ᑥ�XK��sWK3��웲l�����|�6�W�c4�P/�,���5t���woޗ9�ο��8���>�~U,{s��l���F���dO\8�����^oȸ=?���)�"^��k�f��L�'!���>�w]eo�K���N�P\�,���Pl�*;�kɧ�o�l� �}�${�Q���������Ex�s�ayW����u�Ũ������Z�<������1B�����5��|�͵��un�a���-��/��*=�͔�������אּ� ���|#p��Z�*cP�&Cs���/ٯ���3�����#�S�O�eؗ�E��#�t��������	~o�3��33Kj��A/�O��Ͱ�yt���v�8Z�.*�	0Ԉ��Pg�=j�^qd+�x
�n�G�V7:_\�\Z5�%5���O�@�6sh�\�f�nK���P�)Q)`�ۋ���y���x���J�8��t<��\����q}P4���*՚��u-��nH�~�A,��H��E�^�U���I�T����.���_��ӎ��ֺ/���I�=Mn�)7]�LJ��p���������q9�ƨ���?�]�+�j��=(�ê�V\����b&}�;hK��O�s�f�B:L��d0gX����,D'���3M֜?T3�UwTlx8U�� 7��E�8����yTʽZT1禍����[5�[x�f��,�K<7v͋3��)]�)%�U�u��<�B�}����o�o7=t�n��rs��0���^3|_�-���%͈<�>Ѡ^������H�`���e�ʘI��/��^%����R��>��,X����p��1��k5���?�#���ֵ�(���UhL�~�-�z2���a ��4q:����o��9i���ˤ�0��,�ȩMU}��D7(�<�U9�־Fx]w��L��Q2��/]��gf�/�~�6��c֖X�K\�SyQu�B(�yQ�q��t���2UZe��ƿ]��?�Z�WV�Z�e���,�ˣ6[j��bh�d����4W��)�2Q��,�rS|[�P�E��bB��$d*����������s���������Ց����NV}��\��_ّ�"79nZH�B6?h-��nIVݗW�q10_�� �H:�8�h����L_���C���Ӕ�\��wϞ���d�q���UT�������K~�R'�>Ǜ׭9A:;Ƀ�L�����4�`]ꬒ�7�]�v����Ndg�<*Z�-�'�����ּ ~W��f=0���lW$��D���(D��u��SIP���hX�E���IX
�y��6�F���n���;���oH�Y�v���	U���~��D�)�Ut��X����.�Wf�aߜ�p���e�v�{a�}�������GG�u���b�Gl4���)<d8/�}$�V\O��pO�Y���U,�ᨦ�H'�Rp�%1�����~?v���WC�y�3-4���<�v�Ea�ɸ,r\Vҳ��/{8Q��'�0�S��X��k!(�u���?�Yq�v�(s�Ax&���bӹ�B`��r�yK� �� X��R��9R���-���x2��G�B�}�h����<Mil��|:�)P=1�֛�<|ǛeWY/���=��iI?E� ��];�<�ܭ�C����DJ'[����s��K��)�yDoG���L��]Oei�9,7���̪h�7���Ԍ���F�!�C?4���Nd����a�ۏgyZ�aˆ'�˰�����Hu$���˓�0%5-ZH��E�t L����^��U�t1���&7��'7������ݫ�Ϳ�$d)���_2��\"z�l V�iMn����H�.D�:�5sӶ-�Y�� ���\�ы��B�u�*����)��a��V�r�5���1�?!L��)��dFIE��쒑k���ע�!zz������Ul'.f,���N0Cz��` �"����{�T���	'b��C.>�r�΃(}M�7n	6ظ�[����w�<3\goSEc��C��e1yo$��opk7�+�70،��d���>"��3�&k���6�W��o�O'����
�v�k�~�y������`������N��O��%�'�J!�:��;�bMk��Q��m� ӊ���w���ٺ���m��m,<_�ò�.�5������$u�l�T1A��FsoV�؉��\_0=�$���YL)L�2/v��k��g]Ƨ�`ҍ�����w�y���̙���q���ud���O�C��\{C����U�j�}@N�=�t�a11(\����	������ݹ���E��j��:MX����{�ȥ��[�d{*GD�w���%�-)�+�A�^j"(7��y�+!�j��W\���{�U� ��t'��m�2�5�݄��B4}y=�`�up:�a�N��J���U�#�jD�#7)en�6�e+s%�ǫ�}��cQ��Xh�z�S�_M!66�(��8�?1?&=�^�%��/C�7R�\��e�_j���9bZ�1TWP�Ȯ���qV�J�����4܊�AGG��r �k��~�M���ɍ���veko$W�xMH�}ɼu%�o�q��S��ۡu
�����~=j�>��!\L�[S���e(�NX0�^_3���+V��]{T�{׳���Sr�}�QF��C�+�^9 �'(7��1e`YP�W�A��/8��,�`�K G�n��'��ş&<�>�m��߬����M
\h�e�o�H��@h������PK   r}rZר� �* /   images/731a9da8-b9b1-4e67-98b9-c038a7318a47.png�{�_�����atw�0BRDiIiFHw)R"!]"�):J���(������_����a��ǽ�ڽ�\�3�9{cd�EA�D
  (��<2 p{�ĄwW��4�O$�O,� 2ڻ ��
�~�f\�j}a�w�z�Xi-w���˸�9�����Z�H.�ho��]�X�8[-�s>ld�w������~a�'P���e��Ѡ�j���O/=��L.@�;F`�Ĭna�Y ��kIP���U�:1g|F�HԢy�������g��4�]�{��ߋ'H{��F�"y�E��sލ�=�I�FO�*t��_2�/��B�/��B�/��B�/���P���}���,c��$����1F���G�|O��Fԛ�_��o���6-��vP�[�ׁ d�X&O�������.��=���/a����HM�o~�����I�$�b/�?� ����� "� l�B?��A��:�m�Gz�i��F	���q���B�@��ݻa亢T��\G����r����o�	�,�r / �~�?���?�_�r�1�.�f�����U/���^M�9�l�)PÑ��n��0��)1*�7�Q<�����S�o�a[F���ۈ���Y�]�j���^�$-\�P��zK+15�!D���	A%Ϸ��9��ӫV���������<��CV�?��C�.����e�	�O�MX	��_O����\�F���c[2�� ��3���'�� `���§M���-�e!*��]��s�Yz��Wܮ�jxTw̫��=��<�����2�ZI���/�� �2�̬N�PIi����WPߊV=�?M�|P��`յ{�s!f�S� ޭnP��٭��w\+��5t�r�-6��Ep=��tZ�E��'��Ai�t�"iN�V���R���$�$�M{�w@�6P�2�h�o �PW JBV�p�2�V�:&cJ�V�ܹϠ�������O5�W�N'@R'���o��h�I���}-�i?@N�'�!�Ο�G��^�����ר�_T����;g�䑵��U��-����S����w ��uR�7@����ݏ!�I\K�Qz�絜�����T�K��X������'������ޟ��I�v�o���_�ދ�������B��Ĭ��Hp�\�_mn9x�_".g-z#�cddq�s�2:���.1Q�S������.y9�9അMNL�y�fvu8i���C��_�d86����|�=�A��a��ZJ�Y�F�e�]=���#QP����K�F�uj�i߃59C�{��(��椤�y�O��xy1e�t��o��C�G��4�����rrh`Y!���b�l*O���x<d��%?����|�֪ű�JpV&ہ%�=��P�@:rӺn1g��]~���X����</]4I�Y�]��O�����CʌD�Ĕ1�ZQ7�������]W������"9@��j� Yy�%2ec� �,�sJZڎG�P��r��%�!
s\��N��u�M��3etê_�<XP��#��C.옠u<�����l�/2���F�����/�L��������Q���Rփ��4Ϳ�]�r~#��$�z��_{�u,Յ=:�FV���sFVN��V�m��ey�itd���.ФHZ��cA�WYB	�"��O*àb��)�X��;�������$h�5���YV�T��?1)�@��z0�����VEhKi�0:]�� ����MO`nVp}2yƛ��r�tM���P�vㄟ7�*���	�r�i@ig���z�껌�;�u���Y#���]��|y��7��w� �uй.�T�~S���7C��x7.j�n8��٨�,��JG�����������ߟ��kP�|�������'�z?ފu����!V|�)��M��v�UC��1K��8�?i\6����ڽ|��h&]h���2׾}�&��ox{�{�6���O2*��V%9�-|��5���+f?�o�TWc<`�E;�#͉GwZx��e1�����@,wȱ�l��Ľ�c&��৞D&@�挰�`�T�K[��?��y۩������ָyYԅܓ�Xx��{��ش��׸)�9�5<�,�����^n��O�Y�x$�=k�i�7�s�&�$"�wH����|��o�lۇ�Z��g��t���`J�bj��ŅT�:^CC�f�����G���1���R�R�{����W�W�;��):�:���];ٞ�ښ*
�X#��{w�	���&���YMj�C���4��b(�5Ǚ����o�(hm���[/z���
ځ�,o�O{�*j���$�'t����ٚA*r�q���Y���J)k���||�<�F �l}�_�g��v/'��F���i�g<�Aֲ��h
�[�*	�<��]�?g]$����q��(������ݻ� �l[�9�U���뽊˻���}!�%�Ѵ\k�[�C�-���N1�������G����K����?�ZgXcj�`�w�C���@<xP�8��"T�_���Q7�}ify��Щ��!�����f�{6�ξ	�{��
��ԄU���O𸸸�"�>>�g�[���!	�}�����X�t(�;����\'�����_ֱ��W޽���C�~{���E�X��M���T輘��@j���O�X=�V�3�W��C��b�J�ڨ&k�S����C�I�����S���5�Ԅ�Ry�[ʘz��8�s8�gs>=�!�~r�.s���{*�+y�'��7^�nٚ���!�����,s.߾}�����`R"֫�Ñ1��cc���Ld,���J���	X��τ5kF���j}�C�Dw�{F���Ė*���Ɋ'l�(��O���O�Nϖty��;�B�^Ն�	L���?3ߋ���=���݈rss��X�M��R#��!7��
���{ձ�1ޜv,�}[�Z9y�/�8Tˌ D3;��Wւ���*E�;����G�����@'ߣL���r*��-��bT5�����O�(�eʲw�|*X��E,Qu/��~+�{����W������e�[_�+[�V�4�����_[�a��j���vJ~�TPjUWnV���1�g�=]]U�Mu��"�X	��+�`�>�H�z-F�2C5������R��l�0�65��A�B�U](��v��w�=ͧa1`�@���G%� ���IM>���� �5�х�ɪ���О�|�i��@/p��<��/<ǀ�lk�2	"�H�p'����*�5�l�
+��7G����ߞ���]�QQ����)^��>`�hY���s�:��mU�	�;���
�t?l{PL��|<p�w`�K�՛�i��D�/��:�� .�J��ɥM���u�W^��eną�x��{�)yW���H��:���E�c�1���q�\�m�E?���
&8����Oi��Ǣ¨s��:��fFW�+������j�٦?/lʿ8��wwr**N�ޤ�BtY'���.^
8,;�\����bZ���=?����#I����^���@6�@.ه��Zv�/|u�׿1��^$��H$[o���&^�Y����7��7F���48>f�K��b��+av�*�-L+VЮ���c�V��w<OR�_i`�+i�L���v������~!�}8B���f���7��JKV���b�� ��Tf��f�]x7z�_%����@��=Y}�mC�я���7?�T�������uT��x(�ܖ�9��L��~Q��y�N��R���G`ww��?Zqy,uFE�8�3H-bSͯ�A^��8"
j�yA�i΄~M��,N2�}�] ^���i�Q�φ��:@�O�({;���|���fp�+ou,E�L�f�P��F�Ab�'�otźw!���Ǧ1�E.�Y?���<ڡ�2n?v)�r�*ҏ-Qn�N��;u|?*��2'ڊ(�m���؏\�W� �`���\�P�ɺ/�ܜ�'S!lU�C-��}MNtn?�H�HF^i��Ƈ4O�2�.�R�fb��-s1�&.��)b݅j�/@Bwp.]�h�ٻ������B�9��{�<jM�R�^�Ƒ��`2Λ�;.ҝ��ߒ�F/����m/��F�|�:�j��W��A`b��lthH�-sB�2q)e��Ai֐1��O�C��G�b%��&���f�z�8o�H$�3>��بv�H�~�Jytt�w5��4��%�,il�%v8 R"������qQ����ݙ���&��F~�+I�+������HǽK�UD[�3j����6m�X���[�xp]wu�5}~��f���@�:Ǎi���Y����$�X��]l�)�2ϕy-�����̓�U>9]�]�ھi4sp��<H�t�!yu�X[��Y�9y�i:�����riA.�&n��ۖx6663�=[���/����<WTdd��D���Gǭ|2�o��K(�m�6�C�2"����օz���>��WSA}����l����KW>U�s���$���K��ZG���.��������(��'o�|�{ͣm$B�q��!����JcQ����5���X��<S��pvA���#�"�'�a��s[>�C}���꧙��>�hQ�5�OE�)5������jēH+���D�9����?���U>G�]Oc�������6��B���J&�ԯ�9=N5���X*,N8�����Pc��'��o��K�(֑̐������{�����ۉ|0�U����F۴�����]HRY9�'��C^^�:�8V5G�R���s�'u�z&t�K�6О�,B?7�:kl����p��}�QO��U��s����=��е�=�&�LKK����'+�ck��z]N���*H`m�&S���3[�_݅����e�8�7s��VZ�����-���E�R�>N|�[���Yy�GY�6�PnxqsnB��V�Е�}c��Kl�g"�L�/u��ܞ?�u���}�4"����P�nє9cpdL�����o��]0lr����OY	���o7�ow�m�����}�cs5��i�)9G����l�3��κg@���d��J�Ǐ��.���ԉ�^D��"""��FƧ����.��n,J������9�F��WA��>+��<"
��?&F�m����}ܯ�j���N�O�0}.=V��A3Z�^}�9 �&�OI*=En�i����X{��"���?��;F]�E�t������`�d�V+
�}�'�Z�h#1���̈́I��񕅼R|�#�P$[UU%!/�`֝P9�ԬWa*��"�nό9�g����:֘tc�y^ȠD95
�np
g�GqA�,�r�CW+�3�$A����
-��ye�[µz�/~xu�aE�j�[DF�P��8�!�?b� q�f8�򾫫�W����ˁ��-��Ϝ��)+�I�
L��rS�s��"��bg��c�9䭑m��f+�jŽC�#谝-�J�x	8cVf��uCO��Q���θH�u�j�>CՋQ\�"@�tK�drcg+14�	�w"�5��g��V��QW����F�дs����� �ny.@���,���̗���)�Y�� 6���%���nw��S��c�y�`c������[�?�S,�*Ұ�tk�>xTg������W�̆Dg�!b�������ch׫W�4[a����X�T/����)]��'9w��K�o?W��%�"4k���(���2�;Z7&7Õ�α���V/�dS:�B��{����2_�+�#Y�~Yȝ���f{� �;���jЍ�C6 �)p��A� P�а+c�X͐`/���36�_z�*0��g�
<��k��:��P<iii,|+�����i+�Rî�7�zz�n�����SE��($������j'��Ƚ��I��6�����[��4n2�:�/��1�v�����+DB���-g9�mdmQh�7���r>Q�+8�����,=�I)���~9S�&��L�i�f����7"+<E����g���mN3C��"0���.2�u���t����:�+N]iS��_9��=�[,i�,�@��ϵ���0��Y�x�%{;k��oY��jMc�{�6뇧�����1�g���@l^�n�a�R�-�_�@3��>��L�f?���,�2�XSY�c�� ϯC�>04��C������)�nYL��=�U��m�֏���v�\S�@����dN�I5���$�>�D�֞�+�WL,���L����d��@:�c�4�+$�}nO�WN��0�}y��uW,Oi��Ř�'��h��n�������*
rD��?���
o�,�'t��Gƛ�)8i��Z8}�����b=��^ˍ$Ն%����F��tw�ҳ�,�����K�3ͩ5��\ ɢ��ĔJ�PD-5G�>�,"P�1&߹Wбzg�%����������\��lb���(%����*�C��L��$��<�)8�zU���
�G�λw�94�ǒ��h��,Ǒ�ĭGE7�?���q��ý�Y���.N��
`u�g��2L�Jt�W��Hz\�S/��̹,5����� T��ׂI�ς�������>9�̆��؝ט��i4D�n��U��i_{�%K�Oǒ���y���H����_)X�v�.���c]k�o���~dŜ�p3�ΆJ-�)O\�o�Ҙ�H#)����f�8�h���K���a"J'{��B{m��.�m�]�A"�J(�A}�����
e%�p-40'�/V���	�����4����hs��MF����p��j�p'UX�1'�Q�И���f-� ����K�ȫ=̨������V4l�����	���K���Q#NHh{�k���gMI!w������%��މ.k��K2�6p�؞~6ϛW�ȋ6#�C����MHe�j�ȁC����XaMNW������q�9�.���1����!Ÿf���J+�M�(��}�]�+��4q�O��L�]LsR���L���r��0�o�A�٧k�l����<y0��׆�}�K_��_����$^/_��H+Y��^�i-"�8�9��x�����ŷZ}��n	���a��	 ~��.V��ޓ�&=V �Q��x�H@89��>����ԁ�[�Q���Dgt���a�je�O��,�̨�������&�3�_���a���Sz�'�[�¦6����N<z��iLq��Q߷W��@ܞmNȲ����Z����G�MR��������D�!"ΤKN�����{�iE8��b^ܹh'��x���GG����x��O��X�c����p�?�]��f����C�(	ۥ1���렡�	:��s��A�_%+<w��5���Դ�/=<Z�h��~SC8Ź+��������_��S;�i�O���Dg��(�X���&(�(�[}�tW���r��7�	yy�go���b�6��u�sՏ �6l?�W�w�L5�L�	eK()�C�z�:L���!�d���j�2���^�_[���W8���:��+�A"9kia������x�ґ$A�^����ۀ�����]�a���b�:��f.�j\�k�2�i�O0�>�!U����B�^�F�`Nb��j�.�?�͵,�^��x+�N~?�����+b��n�^�z���_�q �����iqf�y����ۡM��h߶�U�(�Dt@� ���Z�4w�t�Vd���\� �K1�f����s���vm			P���cȏ�1�.��	�զ��?�U.��\���짧� �=���]w^�8�~})ݺ[��ys�_�ow4�珻���ڃ�
��u�B&���^����Ԧ�����q���	�w % ������Hҝⷘ�R���U7\�i�3��V�^û���#v����v�Z�)��I��w&���LJ�Xҵ��'^��f,a��yb7<jK��
�˽�^rMBHHX|N�0*ȞO���B��������S2�́f����<dl�	���v8�P�T���Z贚��_¶oVW�d�����1�@�
|NtLH���1Qz���\��Z�SA���=D�Y�`���^���_�]�#Ǒc��s��'��,�0�N�-�z��;d��#ܸ����r醝ϭ�Z�.�W��X��>�}��&�̕����O~�]l�ר���3rϪ��8�F���3�t�����I٩�k����� �ϳr��Ũ���)0�pO��f���Μ���������Af��v&�����]a�Mn$g��N�'�3�:	))cV��尃ޕD
f�1I�ۣ\���T�o��\��� k�7ƙ)�V�4Δ�\` �2�[[O}~�t�Hb
a�Gg�[�Z8jzٻ�߈x�=s�&"K��,�	V�4��F'����y�R�Փ:�+Y2�K&X;�Ov��9O�%�;����,��:�)	M�Ϩ����,���4���V��o��1/!aXCto�{��^�A���ѥmq������ݐ��*&�
)oO#���u�e�'m�E�TN�͑�>�T������&�������¸�Ը&���J�M�X�H��}w�`4��Y�ܸ�����(VI�|n���	_< DX�~��w�,b?���^@\O"l"h��S��9H�����uz�}������BN���������3�k�0�t�b�^�a���L���\�K� 5�F#�Q�X7f�N!����7|7Ѵ����>�C���9�K@���9č6����� ��>�	ޟ�s�<|�N�J�����|����� ��w������m8U�_�D��9�*4r��T���� pxb����Z�|�v�{��x�7�Ή}�:\��J��8Ho�q�<�&��2����P�M����ţޅh$K�sBl�cq����b#X:�[�=ڸ*�߼�]���W��F6�ow<�Ũ	V��m��Ue�˷��f��zw�,-Y�e7�����yc��0::jD'hl~�UD�^�mȀ�='�3����^�d��1  �k��}qd.���^
�o�z��L����8}?��P�;�o@�m��z�x����-�D	�@��M�s�s"w��ŕ�%�TY
��P=��OZ�8��I%!o)$���lN��}�����*{nb��a�|OE���x�� 44��-l��a�'Z��Y �d2�B9{���I$߸�|{���07{�#�OO��#�M�?�GX����JU��2���Č�<#d�����7��:SJ����e��B�wO��W���ю��o7PÌq�����9H�{�:{|�r��-y �L�V�{���fE�~{��o����HԨ��Y;{�7�{�ױ~X6
�P�����d��8W��`�����/)�<I�A�C^���"�~kS�Gd�_��)��#Ω�&�$v�D
��Ø�bE_X�F\?&OO+_���K�`�(���9���=i=��1x���=�?��0o���f��=�r�ӿ�W.v��F>��X�^b07*Xk�?��?���I�|�_S\�.���9VJ�&�!nЫN�W>�-���ݦ1j5�G_��OZ�պSM֫%�䒾~��F<}<p�y%�����U !RO�ŕR�I���*��3,���Kuk��1���>g�x�HFF�IT����8��g@��N�x/^��|jч3�N+��Fj͘SB�na�sfЏ�e{����Q�;~L(�f�2�Oڣ���Zdس^ȭ�ş>6�1ͨ�9U��H<��a�m9e�R�U��v~j]���L5!�D¤�P�Q��w==={?w6]|52n��U2;b��G�݋�/!��Za��0�q�M�dEs��:ꓸ��{佾u.R�B�@&5`�m��@���� �C:��g\o�1j��Ґ��S���:�5�olp�\(p�K?��.EPs��[�n�?k)����=��;@��8p���蘈��`���x����Vt����u��"J�=���t=��>�~�!������U�����Ey#��,?6��%%%����KT{m��X�/4�TJ}@y�`yG�&x5a��L�ҏ��2����l�'stƌ��j:o�k�u*q9A�2��K�����Ѕ�JT9`��4��D�r�hˡ�,F�- 33������ְ���]}=}eIn�I]������������p��/v�l�����^M:/~���,Y$�6�.$�7F�e�Eb��}(J[�7��e�{�>�ķn����Wg{�X���ܠ�W�F��PP#b��ڍH��kU������>�w�|��ћD~U�I���JD��$�S'�2B����;��1�H�v1:)��pqu�R�4������ܳ�V���蘪v&R���
�7p�M��b�~�+˘+�<��X��XvH%���?���>R�kO�o`��MY�ONIɥk"PI���J�{�;"��$�klb�PuV6�v'Dt*�Ԣ���ojl��%�:e,h���8��kt����B������c�Xr��8]�� ���1��_�KI���4*�`"Q��~</���I���˾~,J����a�E:6���|��<y-v�d�n�1��1Q�[G�*H�o4�O�
��?@>
d��ɮ�hcʟt�ɆF�R&�Қ"�Z\�&�"�X`#Kg�uJ_���I>x���Ւ���M��g�;�f(\
!Gt��?���{�d���
X��>�䤈���=?��~UU����{��T���V{�6С�C�V�t�A���u]X��%ې�#`b�j"s	�|
�A�iNsܿ�))��Gʔ<#���98>�Eտĭ5�i[�e!���]L`�=�n�9I����a�o�dJ(x��G�!+�. ����vw������b��ûM*,Gǫ�W�䷅��Z֘�d��c9��:�J�YXXa�	�@K��4x�y%ڬ;�'����*N2M ��4�U���6�Ҍ�X�Eb���hޣ���P:KN�q���� .��ğc�zm�f.�S� ������i�r5�)�gbQ8��S1|�I�9��NX�(#]�һ��VdUZҔ8{������R���t�%�}����)���Mr�`5k���B�O�\�5��:��H�VS��� �@˰(��9�J� �K�	ܭ��o�ȭ$�ٺ�$������Z��EO�ZL$RSfb/1*�N�����G��ZB�@	��g���)>�A����ї�4"���o�v#�9w��TC��w�~\��pO��V�%(,R*�D���x�z���:Hv֧r�U,Y�9�.,�h�)��P��$Zw�4�n_ވ���`iy��dS��h2��=�
?�c�l�����Eh.�UXW�a�햝z1q/���m���E`���w�66˾��׵Ζ�N^��L9`n��!�y��`U�kH�5�nݤ�ݮj~�����'Z.R7Y��9r#�\5p�5 ��8�6�E�K��tE�����B�Ű���E���u��$d1����I��������d*�y8D�t��TW��&?b8ʞ[/�_��úk;=�Gt��R%U�	\H,�𠁓��/��(2��%�s�,�ɀ_��5o#��,�~V58��ZZt��S��#>m#����W����K��NQ]|e�h���e�6U��\��ipǻ�x�q}<y�$E�$	hd(�]��G�DVX��ޑSl���$"�;P���m|?6aڬ�D�cv�Z�tǥ�K�\��ԯ��s�czPЍ���ui��g�9_��mh���"�B����uy�ERM�Y�c� �?U��zDS�˯)�� ��6��7bf��H<7��ppG�q�o���E�i|�ϑ�R����\�⿇�ڳ9ߐtp���ٺ��$I��X���9L�~� �2]������5%�j@g�DN?��>AI/����ƅ��\ݚ�w� Nv
��)�Sk�)�WM@��JF|�l�E֪��|���2q9��� ��OJ�aSy����6,�]`��P�+�'Q!�����ָ^y!HTc��&?���bS�*ꭶUB�u��b,wM.���X���ƛ��%�lN̠��|o`����{���X��`�>3,���ʼA��d��]�aK~���ܛ]��i�~��q��=̇wI�M�i��6�䰨V=�Ez�VI~+�C���š�����n��*�/U}P��X�M"��ÄM��E7��%��xx�9	����}Ũ_�(S�r�9�����-����+����~ CW��߮�Lz֒!��I?���ߴԿlx[ou��X0�a���+��R��D�x��ԣK~��yг�����B_3�I�@?"q�V�w�>g�aɵ�&�]ZG�nɧR<��>|?{�E�zox8])�����xkuVW\R�[J#�ꐕ!r0	���JԾ헓dۢ�{���@��p��B�:��,LC��b�^��.-o�"�K_��vRߓoQ�4&)��n���Q���������� �`���$Ҁ�� �s�s���j��&�$	����p��:�!)�Ztm}(==}ck+1'`�1�@���F����,n�՗0��(}o��YMux?��e� �ڤ�_6�֩L����a��L�äڍa�o01��it6h��Z����Ձ�>�P�u&wz�F[�)eB�z��KP��-ۚ�t�W�:�o��$e;ŉBD,B,�ioz�R�[Xr~��|g���eٴj!~i_���{gF�<�g45�y	�B�cZ�=��t��������<��/h�����,������G��5�Ȳ��A����SB=�7�m��d��(�oO����Ŋ2�94Z���2K�i�٨U���hN'�*�X�#�A��+�p�j�i���/K�G[
|�j�@P'�B�S0�3�}��j1��L>$��-0����Snf��hKc{��ժ���>Qʹw�dB;��k�?��R�+��+~�-�η��n�E7���ge4X���P
��v���Vʘe�a;�^�X�I�=�j���~@���G��������wy7��w��1:�{���Lw���+	��ڶ42Zd�a�0�c$�y���o����0��?my�?C��W'fz���_�33>�;�#~^��YL���b�Z,EӦw�(Xl6�
~��Fs�
p>�'�h���x�rv�R'j=.�
��.r�{*BJ��v:�����\k$j~��Ý��V�R��	�������c[.>�|t����Yg������v0��t
V\O�zSWf�����f�5Udh�����Z��Rf$�u%`X�P��4V��S�Kr�;3��'��lC�C�~65b�RnU����qEbh�{>�ǋ3<�2��J�@7�4�!k�q1/�b�o#Udǁ �@ֶ���@�|�$�F֌�XG����4(�J` ;u��6��wJa�p�l���\Hs������ɉ%,�a�Ғ��b',h��X4T'�	���&UBhT����!XH���@�"6hH�2�&�$IW�ȢJ���8't��kr�M&�J�����a[H_Y�$!}���{H`���S:�m�<�}�5��@ڣR~�]�_Rrw2}rz�ҷy�9θp[��˿�3�lu!8�8`�  nZ�h�q��x�Ɖ�p�X)82�_��b#���S�Ӊ���q���<j�C3a<�u?�4�ئg��aR�M�]Q�z��3ZZ\CD?�"@��؞�R� s3ؒ�|*@����pnf�ĵ�������^������n�A�X�ww4��#�i�(���@�k�O�� h��w
�[e�'�@DT�|��i�ٿ������-���܁f�,^��F,��n��f�l��	D� 5Z��U�3��ٺ�Oސ�wr��_���NcQL���]��]�>��]}��m����G��{�>u9���GZ�����o��T���z�T]h��WM�VP�j�&�#ט&��6s��A(��Eyu�A{�\����ۜK��\�B�����7r�����^�o]O�k�ݔK����	�U}���u�]�nڙ��R �B.���� ����g��V8�-+I�����F�A?����%S*���Fh�'eP	7!r�d�í�z�u��ԉ�=U����VI��SԘQ���JH76�Et��)�}��~A`Sa��g�]�@��7.���vh���t�'t�;�����UƊ�
�6kz��2�����E��Ψ��y�a2�#wܚ�ה-�n�GQX�$a�������H���X��k"تˇ<c��G���� S�r��	_0I���z�1�@ҷ��I�����'!R_2ZB��g�m|%��;���B��/�9K6l�-��ˈ���Ƶb��`���͂mWmb��f��g����B�#�	+�hp��'����I�.a�t)������'��:��6z<�5����ܩmr@� YX�׉���	�n^#g��!���[�0�P6���q��b{�p�Ѓ7z�7��~+k=d�Co��"���-�_t��B�� .t�l�#f�D��&BB�)�xr�qSg�8έ��\9���*����s ��D��
�;��V�
&e����i�S�f0a��0��8�=�ڝ���j�J����ɧ�� �8P�U�~ 6g�_���e��q'Ӻ͍ �����qefjp�Ӿ�%G??΃L�NᜌZ᷿�Z���U츉���s�m�@eGg����+�4��x^��F^�P_~�Q����q�Q�0A�$�h�'Q㶃+�k�M���07�����.x�gk��:`�:Uv��z�p?��U�N�+��J$��Tp��a�Ym�NÒW�qMდW�vݜ�a�]�ӻ�x� ~�}�;g(P��5��0A@۞6<x*�{� >'�.ꐧ/G����/y9BrD�ϊZl1���X��X���t��Z=�GH���t��E�ټڮ���"���~�b��9�2S��#NNN���]bl��z��N��5V"�?�;�9�������|�"9Mk�+�M����U����Ԧ^���̯t�O�+����O�g��O�U9�y{�r@\�g���f0s����7�ݱ���+6	"����./��ZՃrw$���3���\�v��di�L�i��$�<ݖE��H�3��M��08��0�ź���o,�U���r|��`:v��r���vd�K�1�jL"�ΠP��l���m`���X�B>%�XK�]�U�����W������.[ހr '���J�*�־�n���CtD:[4�r��/U'�8{'��G ���O�O�-T���'�����;�}�B��j`P<�;��Ct�=5K����: 7���9k@�T�>gN3�6y�u��q�l�	f�ۈn�6��Nw �:�p�.�H[S�V,x�ר�s�r�Ǿ�!�>m���Q]�:�ǄeL��-��}���#F���:]�,@��q�S�q̀Yk E2��ڞ�B�Ydĸ���IZ�'|
UvI)��.�x�"t5�Ƴ5]�)�E�>K_<U�AkٔE���e���_i���[�	�����g�d�8-�+��u.D�:���e�_�ɰ�Z�k�R�=��za�u��d�p�xc���l�1�V9��L�����[z�����>���g=�:�)墯?F��ׯ,X/���ob���z4*q\�
����v�JV ����8��2���*%�TǍ��ଓ'��ʞc��,-dǟ:�?A�0+�~�~��A���)i�q�����Ŷ0�f��]�v���n�N��db�nV�Ɯ�>/���Jʋ���5���ө��/AUkaM���:���@�D�s�W.׋����lB+�ܢ�Ʞ��A Z�6B(S>Nږ�{*HwR���II�XXƑbW��@�[��/K�rt0A����}�i����"�ji�k��]� [8�P�Wq
N2�\�q�j�k���	�ls���D
�C*�a�6����3+/D��:3���9�)`�9!!!u"��=�̏�L���3Hz�U]A~k�H>Z&o=<��Ӭ��C<�ɳ�t����m�p�s��"�Gve�����N�w
���;#=G����%T;���*gN�U�� ZVZ��/7;{6��.\O�\��,v9뺮W�z�U�[I�Y�lo�&
��b5������w�0��9�յ���σWim4>L}�7W��6�?��f	Z�`P��l�{�j=~L(�{Ҽͪ�.']ٺM@IAI0�PDv�Sq%���	�BѫT�_gJA���n���j�\&L�(�l��6���jj�{%��.~,�:��g6�l�{[�Y�(֧���8�ǐŀҌ��>">P,(���o�7Ə.8*޽'m������yQ��_�+M}x���;,��	�;K<*3
�-��1m��$ ����rt*mo��z�J�
���K���u���`=������ir�5��r�ym��N�Q7em�������y���i�xN��E���yH��5�� z���s����Đ��Ryډ=����rdס��-*���ntvg�X=�[�&��L��1�&�<����"S�NUw䀹�5
�#��
[���e��~s�rNА�A�9g
�G�X	�P�#���^j��
��8:˸�.�ӣ�	�n&�)ݓ��.%�t���t����F#�����K�{�9���s�1,��
+��)E�d����Ƿ%�=�п�S�an�A�=�Ȧ��04����y��lK�h/��g��ld�w��І_-��}@�>esm;֯�zv�m��ph���	_�֝[,#24��&p���骪H�'�8Ο��A+����W4tH@A����q��_���݆nM���-6�]�XU�9���H(�
'�F���8&�6�O�7��6�E��U�@���ɚ�a�Wp0%�8�B�j��=���ef��o����e�o�,C����{o�Mj�O32s#����Ԥ	e~�/r�S������vMB�r4�^\�N�bSS?�~zM�}�:ߪ� �����iD�#�z򶺺�c�s'�U)m�����>�l����?Rv
��5o#�/o��>ؓ*D*�!&&��Cv7	4y��܅��U�mmO��;_��t�D��tv����
b�H�����x{V�y�ΩS<�{
�8.tlݍL0��}h(��,"�V�~:���t=�ԁt����ֶ��Ěkk�w���๢2�Da��o^)�$���xW��o�j�Z�6>4Ԡ��k�tR�d=���Wj�0b��%�y����G�b�?�RΫ�MB��
���{>Rd\}�o�t? ��A��'��]��|hb"^C�(o�����s�m�H0%��n'�G%���9����� �2�gܤ���K��C�Aw޺?wtt��u��^�i+Ǻ�Cp�3L�h��S�a�N����'���	ӻ�M����������<+��%�/����8�� �U����=�l�~�F��{���RlAɬⷵ�s�v�Ew�"G[�`�@%�a��yD	�������Z~l��@�Ra�wBUjd���G.����T�$�<�z��г�l�e"��b��F�����g ��ʧ|���c^��M^ ��r^W�t}�_攎|z?���!91z	��$\^�kdg�O�n슦UzJb߿���e�C-eM<>W�<�;�y��h��ļp����1H�8f'K���+.�2�|���.�2$����W���h�R�W�����ڞf�7��	��<hƠ$��F���x�vF�V���<[��g�yJD��fm$�);Kn�x��gq�3�uIa��V��*-V�\U��lx\'E��&ۛ���̡���y�Ct���`���[Gq7����0ncd5��d��o�`�%@�i���;���T��O�BE��0U��^�����[|r�P��x�v����|�dFN��w�a<d:�%%���)66������:���ry�s^���Dzk����uh�s�V�6�gK�z�y*�����~-��%s*Jmk-�O'�\�W����ط��)a��Hd�f-@����^�.�R�D�߬P���E��qޒ�4{ި�F�2L���ؼ ��?�g�t�l�C:�<� ���9R�#<l�+0��yD(P��H:�	x������<}F�w����� �2�O�,�E����p��Jb����S�\�z#�RD�M7�\}���/�PD=h�>n^?_s�޼{N		����%�n]c�-�/��/����&R��*O9[p+��g�-�9�c8��z{�{۱��:��b������<�oX�YR�2lWp��k�F��:4��lw�ޒꜵ~�fj�X<)@���E:ٍ�I��e�O5yH%~�1f��>Z��ͮ���ny�]
�k�(�(����1#�f��L����$�[4��Y�p����3�pvM��W,���Y���"�5D0Jʄ`�g4�L�-0�+;`� ��JD��r	���&���Cq��p����Y��<0n	�}�Z-�,3"_� N�?��?ƽ�dL��cD 4.1���)I�m�\fN�GNNM��d�Z ��bM ;z |pd҈"��B��z�]D�z���u=�u���9◖�^��@5�WDؙ#��!�>*��d�r�~�� �*/�uTf+W�X"���],��y�rP���pOݏ����7��ُܺ���Y���-b��qc���B����1��V�s��wN�LO-��H{]3����ӗ�/W�s-�s#����;+ոA���d'�ȸ��Z�~�������CK��j�&O]���(���H��I��s[ZY՝>mz�lG;m>�S
y�°2�1E���t�r���9�%<��I�?hSa@ffp�?[�P�a���*�aQ� �t���J���cӎ���=DX��Y����bxZ�P��|k�j�������3��v�}��%�Y�R��f��:1� (��;PӞX��j}Ly?���m>;
V7���IIp#�5�Ubk���ڳ�F�t�"S{_��4_s���)qs���Px`jz���ϩ�8�R�i`�zN��S��DP  ufB<Fn�KX������d����_�4�l&�]���
23�ӷ3�\���u����o�iq�Fstt��1��'�F�b!�DNHzn��vA���yN8�cj0�׽�h�K�-�7h0�dp��f�N'�(��N 3�-����hqH�c�(���]��}eN���-!(���v��w���/�\l'���I�������*�����v��E���e�_y�8D�/.��a�u���^����B�fŤ����y���ا��;�E����!�|mp�y��HLB]�C��8��Z���ŵ��F.����
�*���zW�]ar*]��[��e�e�ۜ�\����״��,#�~�0��8b�����%P��DK��>��,3@|����H�^K8�����<��.(�Eħ��^jk�@_؏ֈ
�nt3&��Vo����&�y�k���yh.�%t,Z��)x��p�����n�7��a��y�>��r�b<�p300�6�@�����UNfX�B�\EdVVV��s���b� ru��F��|�����d�GN����̨��+?�C��H���{^�H�jA�T؂��MH�Ѯ��E)c�W*y.K�e��:.�~��=d��g������ŗv�Z�I�9���QμϠ�7���H�d}i"~U���1���i(@V.A{���Y�c�,Ⱥ�˲�Jm����4y��p}�������Q}^P�:Mcﾉsڸ��{��j�D~긑�I��ӊͶ�K�������2�`��F�١��������~�$�qW��۩��'JX�p�i��=� KK����,\&8'$-�!<O�?� �gnԺ#kW���p@>�u��UB���,����v};ݴ�:�a�ۦ������c��z�8KD77�o{��hl�2�P�%��k��N�^��g���xl��<�,���s��P���W�L�/����ixE=��KUqr������*=gLs�X8�:]C���NR�)�Kȸ`X����T��Mu(RT����`����^/+�n�Ŋ� KS/K�բt����uܮ?�q�W3��O"�����T3���6Ņt��ģ��2��f�'&��)�+)�.:��,��Z���"H������6�͡�Dh\cw��C�;<<�sG�\>������䝟�^U4�֯�<��v9o�H��hW�1��p�=�x;���e��I�:.�Uj-`�p�w6Q��+���;��sT��q����2!`#E�M�øH#��*�L�)��$��d�%%�0���D��¼���#�D:�fA$r�Z���ޤ�z��������T����-���i�+�d�UCħ�Oo����o'"#�X��3�V<���r����\�!$jd����~��w�ѹ">s�`�����p\'q睺�;h�2�x=a��T����t�i럑Ģ[�j1!������]��}[��j~^�>��!��f��;�0�\�X[m��+������W�ħ��5Ж=�U�DS,V-`�Z���I�����U��6�T|��S�����<VERK?��KU.�Ѽ�s>�tߗH^�K}�Y�}A�:�a	�c�60l�gj���j�$hpֲ�~�v=�؁緊�����4���|��]��ww�{e
R�JW��ov�^�N�a��i����[Wg���d�cD�]{B��ʵ*X�q�s!0E)|[jp�����|�l���W���jn~��H�-����a�hW�1���?xw��rV��諓��Vmnl���Z�7���\��D�s3�Ĩu?�0�.֙��o"��0�:J��-����F�2����z�}�l�p��ekWݴ�bJ�6^t�������I��f�uʣ�tKTP��U�|��{'ĶIȞ
������P	���h�©��@}���sU04l����-)mp��܅t۱�]�������������jkk�W3?NLM�Z����Q8����``�`�V�o+h�ͦ��go(�6�؋Lb��ˈ���g�uJ�����R��a�ٙ��V��e5�+(�V�8a[��6ZZ�J�����<%�����ann�W��ϴӤ�_�l�(�f�L�Ɔmb��iU��	a��fǒ� y�\�|se��Jgp&bj*I����h(LJ���T�b�Jd2]�����72����������w� c��������|�X�ϓǱ[����e�� �j���u�O�⃿���-�ژ��B���T��5:4�U/>��;F�JВ3��)�ѧ���x�Ʋ�fBR�A�Kt�-t�%���ie�C��d?,[����-��}�abr�NYs��|���Ʃ�T��~9#n0��(��}rC�F|�����dݬOJJ��Oه��]�����"jh���I��`6~ֿ�6����4�����9^u�0D�:�� �� ��~v��f���2,���V03#}��@���̡�F�^���g���fQ�����bF��nӫ(��gF~vT�+�cW����zfBt�������a��1ii)(�� #�g���[��� zK
�w��;�-����#��x07�H*��4�^|XfS�Ħ�S���gג�$�����ش$�5;�F_^�P�zbVk#&''��=8_QQ�7�}��#]C���6\����"�~4%�w�3_�ň,~�N��<w�r|=tX��!ί�cÓ�x�:�i���U�������u�&�1.��[Ϗ�������'�\�Hb�P'�fK��E�Z2r-��uP���&_�'�L0���]�A�P�]��|�V#���g��e�'`�9ȹUk�Ϯ1	}l���1��=%9�z��i�:���Zofͨ���:��fbb2�:k�4�� I�c�È����}�0x9�����H'kfc6�j/��[=XR�7p<o����/�ר$��*X5��p�~	�py�R�KϚ,�e�~@�/�<R� ��C���ib�:�%�:�El��y���k7&�u����ՠa��w��O����*y��{{�{��%!\h�1�l�X:"Un��-����)�D��n�s2rB!~�M�y��>`�B� _K�y^�V���ܟRQ�C�,�-ٚ�N�Z��z���4,.��*o�;����.lH�X��D:��q!Ou_ ��"=�������v���L��B]�;��4lN�#��K��z�����u���<+�V���8�v�ס=���F�>A&)�>�J�V�G&Y��lǘ�k"�ˏ�3_���vl�v~�q�Ȏ�����ZZJ@�Y����&m�:AN��qz�tKZ�|�f���K�X������ԯ�͔��H!�����{q@S	#,�rKHd��h��G��c�I�f�2��Dc���µ�rO�rWnX�����Xv��fb!�7�/7�'�r1Ow�z[`ߛ/����~�����r-D��� �8�.?S �����$>N��RYG|٥O�yo�`"6Ɛ� �5q��R����]8�?�.��i��VZ��wD��J*� WW�����Yw��E�NA����y���{8�q#�N��ɛڏ�)�����f��,3��-��~�>b�]�|�x�2}C�:nvX���kCi�X�3��7�i��"�i\ 	��:C.,i��*	���2 s�j(nC�[����E]B �f�|F~���P���ɤ����˗����
Ģ�b/F�q@��<�36��J�yPh��D����ז	u��0�ÕR��k�4>��a�EH���L@d9�T7#7�wc3�F1��';{�$�7)iu����Ք������h�Bޤ������5E���ܑ��6/S)�v7X����>�>-ȹj����B\�jC��u��?!��K��:�j�J3r��: y~b��˜p=�|�JE����BUz�g�m?�7��4*����:33s��y�o[�(�<��oYu�h���9as�����^�j�,��͝�\C�h��X&T\�1y�)U�~a~������˱�zF�c}.�m?$\ܙ�5�7t��w�������T�3YC,r�@��h����5#�?���#���V�kb|�
���4���+�G,Sͷ|��X,_-O�L�51j�:��_�rx��x	�Ȟ4��z9���k\w �2�2G�g�m.���g��-i��k��i�Xz4���u�U�	Y��B,#x��~{���@~�9����;ޞk�'e\��k�D�b�͓Jef����	��΋���@�L�C،�)�2E{�����@�����ڠ��ƫ��P�x,��X�⹎ZYu�)���u�7����)�ΦN<V�"4
�]&�������LH���B8�"��ѥ
kO>�jɻ��Yt5�:E�J������i^�hޜ��K;�O��3�EZ�/"�:|������bZA�-*�j>G)vK��.&��/��J@:C����}1�ٶ�-���N����/ӢӍ�;a�	�%�]��[��N0�\��2�������K,�b0�+�܀|���N����u�&nu���,�Y��|��@� �6ɞ,%�L�[��	��h?zǶd��GXZV�I�5�$����B�N0���_Z�_�TU�����R�a��z�Tk�m��軵�\��*Ԏ͸j�OZ� �Xng:
$1�@}VZ-xת`@G��+�j�E��C��u/��4�����������O)��N����&� �X�7���૟&�f8���F��=���.
<��;��<2P�=E��u	���b�� F1Ί�8��;�Y.+��z�B���6%�����u9r�W��
xt��Hy�3W&��?��i�jn9�ߦAR�����F���w?�C_�Z�g��$���H J��o}�����O>o�!gk������2�Ç#�L�^sv՗=�8;�N�q��f�		0�z�X��;���m\���bii'����G9������[Z�Lo���Q�'�ٔo��N��7��м7�vl"�=]�tCՕT��CiC��	瘑\��q\&���/ڗ��a`��j�nۤ�4g �i�:^?c/p���g�2Ht����KMI�����q��mR��Ǉ���S��L;?W�fS�'�/�ј�q�V��+ϡ��߲L�s��<R�`���̩�I%�]�2�c����y�pA`�\i�8�h��Ξ@AA�����0�f�lѲ��Hb�Ԡ�+-+����0�z��E�NP	7c���Iם����ɺį3vxh�b�$���\Xe�L�_��R���]]�<��e}�
�8�Sg�U�[�I��V�U}�?��z��!�����7}1��w��k�{;�;����3X���2�P�%�_1dK�$?A������~F���ф L��wm<7������L4D_V����ȅ�zt����"i���w�4u����3�	�V�WZ�k^L�[ �#Br�.��.ڄ���7D���VQ�Mv��Go�����Z�y&%eU�x��ڙ��w�$�f���?����GG��Wj�~����~Ziv�{.W-Zt4�&EDD�d-9q]�/��6;�P��t�R��cfZ�ıh���BO�<X^Tv�J0�L��<�{ʢ�v�H���SV���N����auf�Z�}&�!����i�̄�G����3�����I��#�Y�!~d��v|�7-.D��H�p.Yfl<��_�'Ët��aJ���.���̛R&��P�Л������ΣP�=��;ڟ���zKz �ė�i'��R`��F~A��CX�<AT��R��:}~ @O�`
k��o�r5�!W�'xc��ɦʷ���mL�o��H��R9���hx���PƑXzְ�� ÷j5�.w-�uj��+`��c��Py�xMB����u����	"�4��׭g�뵍Z��J�2��D���S��_���������sz���l�׵��߀<�R
�9M�*�4��]������ �W`=ۧ^v��@js�u�^?֎_���R��\��%��n}iN; �������+_���{[<�ZV��s����7c08�4q��������Î��3�>'���0��t���nZ���p����`fjZ�2V�"[FE�Yz3� �8:b><��TP�R�j�˴i����L2�oJb�0dI���a33 ^�ņ����x�H�۩�z�L.D0�w����uP%*��\�0B��`KP�iyi�<lB����y�KM<���ZԵ��|7���!��*�;�)�{��-�:>�$=�	��G�A:.��X��H�pc��g����f]�89�,9iBRl 4ÿ}QɪfB�@ ݗ�t�k|h4`G�[:[�i���q~}~�v`а���I�c�e_�Y���Plv yz.��~�p&��	���K���׶�ܤ�;]À|6��ckW;�)�/6��f��5 KO&(��L�v��>Kj4Z�y���	�p��)�7�����J7����d�J�L���TW�m�d�3�",��~�z�j�.S`]o������\��ӭ��r٭�gu-���ҍ��$���̄#�%�os�I(t��p�GK~�̴���]���?	v�buӳ�1|?&�6:PN��Ƞ6���:-yG��ܑ%%��;=!��qC`�|1�#$x�ᜬY}�h|X�p��t4�_�����k��0�dvX=t��X����mV8k�[J!�PXH�[�&U�8��f`�`��o��I���S�=��3,�"����^�7�\���`%�(T���'&�o�ҭ�޻]w�;� t&�����0��Z4� �;]���.�kjm�kS�f`�C�OH��B�k�h���|��(=~�.�����}�E×�4���#�	;0���X�KEb�����`�+���Cq�9OF������씵����.�:\כ!���l������x!$u����E����ln�3��x5�?���%v��'�ۢ�mv5Q������N�h��m3�[�1	��@ڬ��?�Hu.
T�!�ku
�1�&2}ϔ�g��u^eۃ�D�NM�0�S}@��ėO��ߪ�Ҩ����w�JTh8i�g3�(�k&�fi�0�aL����v��?ae���	�H]V���t�=�qX��@���h�H�"	c��P�j�Ff��:%-�a�R�`2?]/���N^p!��?@�UY>$��(\T\���瀳];Ǳ��>�B���V�j̴���zI	���r�����LW����+�%����\~u�֡S�,�nX�M+��=ۥyم!B���}�o���p�iĢW3۶��&�T�|*�dҩ�[������rם_��Qf8�N
���3�G����[d�6ĝ�*���B���8bFO}JB���gWm�\&��a�K�aIz�5�\��K!J��v���d��k�k]8���G���"�2���o�#����+)�1��������#�Y\��V����1����'I2�D�Q5�h�d�3���5�Ĕ��i�[H�1e{�[��e�s�j_�\K@"�����]��J(��/���VlQt�c�1I$J���\z�_�ߪ�]V�����>���yd+աl��լ��wt-�>d��&-�}�ĉ��|��<�l�EDa�kgsl��i5ҿD,�Y2e��h�`z���t�Rs���O�9��b֚W�Nd:L�C-M9�Ro�$A�D0���#6�6sB�\k��������'��hdjB���?%֜G��L�!æ�E�MSI%1�� ���j��w�I|\͎���;�+>��qBOO���2�i#����0���{��h��Y�o0��pf;��oy$A9LZ���R��P�H�vc#����+��L���%9x��j���?�#	��&�Y�0��~��*(x 1V��$L��xdZ$�;c���V�����Ҥ2;i�z>�c����\(A��(� z̉fӼ�P˲R���f�"0�Ϧ1���?<�\i ���G��
lNc_sn��&N�ʥ��W�(��u���:Y��4~�j�i�s.�L�nT��yf����s�9Kv��t��m
pl�X�� �U���3�qx���j��H����V��vp!�kIƎ������ a�#��������ۍM�q�򯥥D�2�=	C�c�$*��W{��(��|�V�/"Ô�D��3P�#���0�l�X��}~�\��_��u�D���5��W�(��*���S�:��t�~���O(e�]{�vAWm�G��<97�)����,ܥ���������-њ�����uF�]��8��I,��;/2,,��S����`�c����HSH�N��˿'�Qw������UB��+@9%���B��������ey�#���F�Q �d:��y�!�IEM�Ⱥ�)v)EpLC�?��5a�ͷ�\��Q�O�nSvM�H��/�|�j,Du���
%�uuܰtظƮ������(�f"9VOmC���Kӥ�硞[3CgG�xM6�E:^���v�.~���8��uӬ�������d_�D�P����4�]Vk�>��`#]�����߃,Uӓ��@3|�>b�~�.kw,7y�V2�|cKL��σ���� ='>����)�^+�*�4{�V%��
D�%�P �i<��C*-Yݙ�� 5;��/7����U.�>XZ�4�{�����@&%#qhS�����N�ޮ)f$s>5��1��'��Kz]k낟��=��R�R������'h�`HTʘ�ՙƾ.[4+Ѱ:�Jf���T;r�aS|�,$�q�}��~��(2�\��dQ���v~�jjZ�����y����,��_�7(MOwm'�U>q�>
B���kT�f����c�cs��'������IAV�(Ə�A{����/��nw��9��5P~�'Fu�)���m��-e��r��4���3#0�ù�]�dn��%N���.0MR�����T(���qF2�}.=aW����y�e��n*J�a� ���V{�V�:e^��jo�V8JTف���;���j?���h��/�!�>��B0IJc�m�@��-��>[����1	�N\4R~����?�Ou�'��Q6�+(���|����Wf6�Y>�NC��;gC��2�_Q a�^zE: ��r�U^a��&t�Ɲ�BT�Qll��|�]�OJG;3�~O����o7(���_���YA$A���j;����X(�ҝ�V���N�.{��12��J�J���w%�~�A�����+����D~PQn��Q���������a<�W�?�m��f���$�_�9u����H�[�T]0-�o�'B��m�m�Q���Lى-�k��چ95)]��-p���" �%���Y�Zȸ'G�hC2#�u��`nU��3�'�N�I�3+q��FU�M�f����3.//o�������a��#�������M���%��<�[�yl:���v+��'��SK�/P l5�bkN�C���|EeVÕ������u�\��j@�7�`��8]*ܲ������91�D'G(�LϬd*�ͦ��3�HK8P1т�����dL�4�x�ì���"�xZpqf AK��$��&F��Xrl�wF�2�(�Q��V��eWR�ܷ��Oc��,TRݰ~�}���0Ϋ3�i�%b�xg���w����D�z���U�.l���c��B�c�� d�<���&c|3x��`����M9#�ŲB�0�V�{���G��P�vD��#��J�@3%sɬ# ��t$:�Z��jd�������_#"�ccci���ge��E/��: M��H��ڴ��xr�>:�0�[-�O�v���
�yB+�w���M�7_:7!�h2i����쏣��u�ѝ�WL(W�C���yf��������GT�(!>]�FIb����kY����N���ω�LSLu�sф�q�⇯�B�~�ȇ�r��5��^�ُ�_�)㕐eM��m��}i��eO>y��<�r��8�`tպA�J�������?�-P���	�$���t�B__�5�"��J���rԑ��{������j���j҅Zܬ<a:u��_�"G5�?�/���$���3�� @L��y�I^�I����S0c�0{ވ�D�L7������P�/"t�I�?jXH�ql��o�uG��Pf�$�_��V#�E�mj���}+,���P2�q��ˋMfQ⵶�m�;���8�,����0.[�o ��/����gE�P��7C�_v��n�����8�g掖��9�+k���v�D�p�lsU�CC2%>ݩ|��[>X�<����|Y���>O<��W��ܻ�@x�t�uL������>��j
���1�A�>�p>���)�g�y����c֒P�Lb	��[��ƹ�be�}<��\��[x~T[�~J��COF�ܸ��G���0�\�Wk�oɄf��ZA���υ�����P��A1�I�8�e�-+2�l��+�7�S��_ O;�mM�u-RC+����_4����8
��+�����dCEm MKJ��f��ˆvP|5�����Y�%�``��5EԜ���ʵkFz�-;D�S���)��we��B�?��C�K%#|�8�������yS�z��ǜPʥ�^�
�m���
��yz)�7 !c=���e���2��'�:A�C�����$Ÿ�N���Wn{�[�2;9���E�uKM^���Q#ý6W���o%.i)�}`�U���)�����g�_�_���ov�>'��y=����˗T�v_ ��}$6��P\�s���� ��c��A����b��(g���'�U
�Q5���Ӱ��� ���R� |3}��,�qS�+@�P74���dS�����u�rw��1}��4���uyR;�r���N �������s���c���%�y3�G���&��pۆ�lks��p���!^侍���8#��Y�?�+d��/����4T�U1+2�#I�寙ѿ��;�5�W�B;;E+�v�֛�y���M[U�w�5ی�X�P7 32 +2F_~��Ź}���}�n����!�;����I;Z�	p��JIb��=����Cq�ɂ����	/+	O��"�o�m�wO��eⱚ���p�W׫�T���M"�q��t�[�8��2���jN�*���.�"w��2�[��Oı^sI �
5z�[�:4u�s�Z(1�����_���	h��K�[��?ihv ��G� �o�L������ְ����rP��25󣀟]NN����)�����E��G8x�Z"؆<li0`W��? ���"oi�<�K��+蜬���"q߷��ї�p
V�x�WT����!a,|�˫N���b(�U'��1|�$���e�Fk�z��<ozB�2��ǩ0�l����&H���1����u�>��&���BM^����1�/����R�?�y���8f�>��ou�x�_��dxs>�ޢ�w��L�(A�n�٨���d ��Hܬ��,�.\��M�:�؁�c�(B���qJW���t��}9L�_��������s�6}�e;���0�O�t�i�oSA���P!��S�53���/V������[@�w�!|�r[����A��=�m��P8�����/+�@cj��?�e������	ۤUY�-HN���΁��� �
(T]�7��"���!��G!�R�-��h�?��!��u�L�C����M3�����Y�'�x8�~5�w���	d62�+m�$N��/�BH��[���Xi�}��{V���>E�d��`Q��6GצV_�lߪ��� Sb�N[���?ȑ�iil`�`��>ԈR�@4�_n���U�w�������A�H��z3U<PK��A}��9�(��� �dRQE����a�s���X��M�->J�\2L�[ǭ,:\Q#E�mr��N�ʔ$ݡ��:Ŗ�;QW@k�d,�������3=�m������8_���;��'��z��#"L��Ko|�N;1�(N������zV��wD��36�SN���{�l�̹t7�~�y�3��,��r�]�N⧊_{�.Fa-���O�9�A?�Az�8>��:�qq������2�bt����^|�dXQ�q(���B[�[���(�	U�Q��͠^��.$�$7RL��]���6o�W}$�?�K�5qcc	:�x����1����P���t2e�ͽ�@�����J%+��h&���w���y�SQS/�ĺ�z�!xL�|��
Q��\i����Q_�<�6 i���*-3S�
Dх�?�S���gW�����]vI}�����,!|�����������W�_��|^���&Dm��f���?>�8uz�ܞ��$%?�EEE�6��9�7��KѾ���d"c�jO,�2������~Lg3R����� zL�����>���ڟ�����N�E��ś�!�^n�_ܜ�۾�,೫�ܻ�c�!��/-�x��g�D[Z!����Q�6]��_��h2����c�}��ޏg-a[GS>�JyX��N����h��eQ'����U�zH���C��+٩M�2֭7m�zZL])\��(�t���[}��H�ۿr�V}�0����ŚW�j�.y��x�'jIp;[� �:�J�U�`�	�wk�n��x��8���l��f=�Q��ކmr������-��O�<|!#�fe3�My���\��>��q=�B�fX��Pe!�����}<4.� ��T���y}w/�Y,rQ�e(���&O�1������nid�jrb��ҧh�q�p�'*�R�ZMH1f1�J����e7�G+!y����=;��a=c���yn�sJ���,��[c�U�1sz1���e�%3�Mg�#h��Ӂ�s^M�ǹ�^�E9C̠��j�������t#�b�P�wk�\�_����i��밠#��h�#�1��F�Z�y�]�X��]�׬���6}딱����(>x�ÿj1�}��ȰQB�pE/FM��$��$���b4�l�4���(��A#E�!��9dEV��}�������Z���Y���y0t"*�Ad�^�=/S2���Yl�<E0��
���K&�Pc�i�&����	A��+�����G��	T��Fho<��.�'�A��Uǿ���>�*�0&�3*/�:?�-q���}���P�hwI~E������[o�� J>�ek��G�ϣx�;�1���s�	���*I��� ��}��K�T+B��4��#%��>`���ϣ�<�$��bu�	r�_��_�k�#0��Aԥ��~�X9\�ܼ:�I�$���;�y��~�82�f?zq��c>~���|i��n�fщ�'slg�sO4����g*Weq�U����Z�{���W���Nw�A P��y���/'��X�C[
��'m�P�X;e���)�M��{��.&��y�b�sl�/�0J�k�}��d鋈a#ƈ$�"�E����h*���RŪ=���"�T$�H�d�&{n_��1^�1S����YU�@�9�qJȽrp��s=��b4�W�����J�Y�К;[�-����F��Ǳ��C�:�˗�;r���u�C<��|���;r}UH���kP�]���l���M��f��y��)t	��/=���y��2�YZ�}7�ϳs� ��M�㌐e����r�a�\��}�H�����.�&��zn���ɇ_����2�U����v�}�B�6M7��Y=;W�sRb�����#�3�Jc�Sg�r0 �=sK��q��S<���[����/���_�~����|�������������+�a���i�k1�8yO�]١�l�}�1S��I�MJK4Be��V�}�RG`�_������-cA<�垆����g%[~U :ߚ
Dn=� �p���;C��T"_2�A��"�{�VdTyvqs�+`c�/��Ϊ�@��uF�$Q	հ�:��?)N�1ja���#bC��eg�L�p�%�c`q�Retĳ�S=�k�$(�k��nm�5Т�rc��X���Ҁ���J�_~j��Y�y��>&�F���+ KY�Y}����;�[�G�z1aeQ���6��ʕ~W��i���j�o�z�_���xǿ�J���z����1I8w�n(��0�AZ��+�Ɯs���&J�D>����+���n���C�n�7;��:*���o��/Y�~������)��+ul����@E���3d�~n �H!{P)�AA��<%�/UU1��Zw�B��f"���$ayS%�3^}�U�կ��w�\����ں�y��0�}���������|1��1��F+E�jr*��PТt�7�<U1I�2�Y]��*����bC�$�4P�hxt-������H.�B�t��q2?A��d���"�4S�����$�yP���ì�e��FawcMG�Jp��H��f����~5���&-�j�V!�/��a+��,����,ڪFz8�<�Ο���H�	k�����	K�Y�Ǘl$���T-�[2�~���n�O��*:N��.[U��cO�N�]��������E��L�vN6�HzI�%��u���s�:���{B*�0�-��.Т���+�i�t݀�����3�J)E�t�"f�����;A���]gl1��vp��E뽧���k�!B����f8�w�vh�Q�%RJ�|�I�_������ʫ�`6��裏FÞKܺu��(�����w�3�N:Y�t�}����K��0����P�\h]pAK��\T0Н��16��le�� i�岃\�k)P]u\�0F��8����d<!�3t�#�-ٱ����<s�K	)Ȳ�#-7M�d2���t�h�4�咭�-��`4qtx
!1Q.��;w���X.�Hl���/��O~���W��-�����	�)�������s9���t�'�ʠ[���4�Xgɢ�Wh#����Jk����GH=R���$������+e%���v��hb wN��5�j����X&�At�z�2�/[��YM�R�IC�O�U2�{��*���B׮�9WH|#��:�{d�����`Z�0axOa#mk�6p~|�o�AUU\�r�Gy�W_�:B����T�L޻Y�k#��a-x��H达2���jI�#�v���=��"뮻s����r}�'����dw3I��Q��������R���N�}� B��n9�1���Q��������_�	Y�^:qw��*�_O�΂QlV;�m�
�}�1K�E��Ӑ����Dd-�g'���W����k�8-��B�Tx�lL��=���������"t#Uy7!?u]�\.�)��[|���|nOg��Xg˓9���x�y�fGLM��;��4�A唐�� tc}:~)�bݮ�@ڒԵ��v��"헵6`u#< ��.I�z�T�`Y�WU��,�4��=v�z?�*o�(tܐX�H���A�����%â�_�M�M,��I蔖UX����O����.\ؙ���>��x��>@�:��G!�����'3�at�9<<��u�QpF�΢U�ё"h�fR�d2��k$@��Y�i�tR��nkT�@6M�R:8� ��!��YEH@�Ep��"`�ˠu�av����!�s�Ǣ%F�5�'oE1�\����>�Bz��2Xǭ�7p��nB�|*g�����Z⽡(
�AF�Td�$�5G���L&#�A�њ!<��px'B�$2x������	<0b���#k������G�����<���{7�x��s|x������N��Y�Jb ��߅�>�]�MH��2��'{�RoVq1�Z���jc:y�<�i�-%��8��X��A�!�:�m�N���O)F�BI�Hr�RuNYM�x���ܭ�ΒK��D�ED��t��I����퇔�1�G�&�E�7MCk���:���RvQ[6|V&5uӄ{=�g����T��>$�"-j��YpͽEK"\::��dY���<<�!1�2V��U%խ%��`i�)�M���������l��,CuUJ�p><��vf�t���6�i:0�>�m�j��A6�S�A9�
X�Mk�������(������u�F�oV0��(e�bQ�XT���Z�3$��dL�V�4����z��� .8���ReH�k�?�ϊ�@[սwS�l����T��U�������bq�mՒ��ԁR6H��ˆŢd��gkk��������tK����t'���4�X��t��=�#$H�Ur���n���80�R0_.�� E$kC�6�m�|�`0"�%�R��,�#�"t�4'�.\������,-H��������|�0��a�� �������'����eYv�+����0�/���6�V�Tj�:TbG�fw°�8�%�Hc.VL�V�v�6?�E&���H��j%���c+���}��ZՑ��ۛq7���0��h"|tU��bh��ӆNk7nT�6��z/�R�_bf��&T����lmS�%��_�E1Ⱥd�����u��4!��li���*��㔽J�1�z����3���"k,E�#�vnJ䊢`4u�d,!D`U[��m2Bm���*�M��d�����Ywv�o��ꞑD�Y;g�b�s���Y:�H �I�l@�ò��˪YO\IUQ�q-BD{n��qqf���ҊLed}f����c-m�TU���@�k�,U�.�`uY�X.���oR�D��Lt��9p�{.�HdW]Bt�Z:v�D�4F�'c��Q��gq�*��J�;U��1d:�W]Tkh�&�N�	���'�Bö���J��m<��*�lh�`0`8�b7͘��ֺ��,��>*������fT�5�e��z0Y�(��ô���y��zs�����c��W�:�^�x/��k�#�v5�lF�5MHҕ� r�NU�
�5�i��1�咺���w����������^��	�@	yxx����˺�)�%.\ �lr�T�X,}�+k�p[��n�;,��Txk1M�G�yTdܧJ�fu,���^b�h�0��*)��*��l�4r�"Dk��r��W:��g'�m����KL�#L�Zfg�]�s6~s�~�d���� �ǉ;uY� ���a2�F�rp�Z�n:w���j)sw�TgXo��n��a	�n��Ȥ@T�5�^4�t�!J10�L&�Y�[�Vz����4-&��:��.�������M��kr/�]���;lkY֑i1�!u��Α��<ҹ����@H.R^
I4�[�"���AeB�-I��Y�82T�	z�*�.���ߺ�O�bGg�z7M�q��<�����B������������������O�o��C�ߤ�+�8��!Sj� �R��D�g���S	�Vk��Y�
!Fd��Ak���}	ӝ��U�cίT�H
��*�OU�x��Z�����l��O;��Q�=M4��?�84͝��:�k�$���"%�I�fm���:U�u$�:�΁u��xL���jג�Н��H��������f�X�MP�6߄�eY��y��spp������~�������'���a������|����v㽏��2�_|��똿��g���*$wrK��ևU�V�<�tfS��N�D���*���&U���|
����4���UŨ���'�{�t7'�;E۶��*�6�^�f�Al�\�[��.�.�nMZ(�"$I�(r��`8v�Z�ؾO����7ϋ��V��X��-�gd�d0�G#��>Gl�'x�p��!��NuYdvƣ����oz�1��mM��XS��+4����m]��H{���r�+��#X��T��P��ϲYuC��jZ�3�u��M&���m�3,Ok	�p0 �xe����K�H%T�._���mk�m�ٸq�F�d�M۩@��~2�E�c�kR���!�8��T-M��R	2dߤV]�-$��d��"���v��;�D��vW^���B���ɻ��J��ܙ�g>�a���D�S����.��D�l�$P*���U�7�5��B:%�)�G�����jVhwv���	����&;wV���Ա��E4ąB$��;_w��qbU����Bk�ai�M��2(D�UL� 72Ɛe���b)q4R8:p�-BmV$5K��{w��Q����b�%�_{�G˲����=����=�0���|��[o�5�H�U�R�ۻL�v�ƀ�ij@a��;��`ɚvT�B����I!o#��tՌ�"��uLTB�Μ���`m�&JV�mUS-�Y�1m��8���3�Q1��ѕ6��\gq0JJ*s�9�I)ѱ�,\`����)��yz+~�"z�󂶮OU�֫
��#�w��ݯ�m���U,#�W�s�| \�F�(�n�:g����%�>��ј��}��2h���Q��p݅��d�T���)1��7���wAH��,#��!��k[�<��"Be��䘭���i��L�Y�J���8�i�s�5Q`>𢋞�I�*�G��-����f' S�cr;�άn�x^<��'쳁r�"�x��3%d��{��%���v��\�z��l�s��Lg3.]��L�����-�,�,���LU�m(�%y��4M���u]3�ϩ��7^{���#nݺ�����nstt���1�k1uKkB�n40�B*��K�M[Q�H��@ T^�A��J����^�&������'��t�H�䴀Tx�J|7���I�/-䜳���β�5�o��B^���<�@w%%͆�L���@�X��JX7��c��[G������W������tl���^)T,r(��>,�Øб�t�*t鐸6�y�mmc��a�,-L&TČ{�iM0���:tnb�X� *7MӐ��ٖ>>��甀ݭLĨ��1�ɔ����:�Әv�w����,��rLݢ��m-B(��Y��X�Je���5o���S�ɳ�S��W���F<Lx�H���o/�)���0��M���UŔQ� a��Y��-���:�ll�(u��GY�����|kZ�p�b�3��8�:�R��������~"H�EH���\�6��X��~�A~�m[Ο?OUU�6B�7h��UY49��9�d�n��*�U��t_e�����22�֞yQ�Y6`8�gy ��8�&�EH����d�Ywj�Ɋ ;�Պ����MEۆI<Uլs�H~�P��LIb�ͯS�6p���%�RO�{��,�*T���ȃI����L1�N9�{��t��O?�l6���sLf�L�f�z;(�t����*�c��9�+�<$F�Rxf�A��ڶ-^I���t�B�ēOv�����b���7�q����n���w���`?$^`[�a^��W��C�ض� t	j�C�5Ut{I^C�J��>¹�O6�_5� b}Ә��K"�eQww�N��s�g��H��D��Y�S��T�t%B���$#��L\R$#��\Y$� ƣ�
��D��[2u�\��\�v��D�?�Gf$z�1�9Y��S�KNN���=��;��i�J�]g-YȒiA��b��H���d�-~ҹO������"}$�F��Jb�����b�����k���o���������~�K�0�}0C4M��GGGb0�};�J&�=m"�{�K� �T�_ۑj�8��U�ڝB���6X!DgGܶu�#��J�4�4;!;�����ݒ�����U1YN2[���nw�4�&m��P�u\��,"�I�E�![[[Qsy���>���~�� %B�y����I/V��䮝���&�De�$�����-��a<�?�����������᰻nm�>�G�������n��]]�knj�l�[��j	1�2 F�)ߴމ^o�Xivɬ�b+K�6{99����]Ƴ)�=�$��^�駟�����s�,���:l���Cl����Hn�SY��,�CMkP�vM���ޚ��ɀu�YA6�u\�����k<߶,NNN�y�:�{|�_��`��7oPU��&I����&`�C��~7K�u����`�j�r��m����[����P^�&�'#\�p���p�8��6,N: zT��+�4�i�R���F֭t�7CȠ��<5.��k��mJ���`2�`ZC#<������I�{Up�&D�,�܊�|� !Y�bmN :�����x�>��Gfr?�R�;�1ݜ�\:��`�H�{?�sB�C	��Lk��b2�ȳ<�6�-O�携�������#^�������?��x��>`Ὃ�^su�X2�QZ3-�0�T5�1��k
ŝ���	�a��>$gE��
�Smk:�rӶ������%�On�����Ƿ�;+ )�M�}�Z����}���ॻ�3�g}N:������-&��)��J���ƍ<��3�?��.r����_JѴm��^߿�K%fw�M�}I���5� ӌ�!a���e�OaRR��`4�g�X`�a>�3��Fkѐ�ƊxL�L�oc�i����Ϯ�һj�6�OWx�*׽�s��"���*��EY�ላ/r��#<����9w��W���{���,T����L��S
�D�
A$g��"��S��F�2b�9�E7IKT�t��R� +��,�zZ�BӒe��|�,�]�ąK����5�'>��Oqp�&o��o��&�x�\�]�_c[�i�
��BU�G�1�d� �@�s}6��Aʄ�^�6��o7~���M
N"�G���V2���
���|Nۆ$L�,&Ŋ�zB�����J)N����д�)'��8����k�	]��j��c�6UW6�6�Ü���2>� TٝsA� r4�Z�&��~�D�}��!�dr"e����"���X�P�ߧJy2���Z!��ŌU�?[��C��Eq��{3��y�S��%�����	��[o�=�2&�XF�o��V����կ��G2����m��abu�u`#+[H2��8^��8UU2�<���p��[T��
V��6�\�L3OhM�|1���ocj�H8)�6�Bx�]2�#v3�gd���Y�����6(�B^����oLlN��~T��U�յ��`0���5b[��;����i�1(��p�<�	82��ӫTp���N8��7�P�ޔ��W�5��$$��GGG]�%�;;3`Ɵ|���d�Ԛ�Y�V$_mX3��a��D���1iK���Y��%3&�)ӭ-�a6�Q6.�Be�e O6�h��d�ǁ㱽���۝�l6��*��)�]�(��I:�X�6`����2�v��T!2.� zA ,[�{Y<̤hᝣ1-R(�a�<�d8�����6O>�4��������.Zh] ��ڟ/+d����4-�9|�M!�bD�r,2ܫ����b���[z�O�~kQd���x�L�L�R��68{i�d:�6a2���&V1���a��y�_��K?�Qn޼��7x��7�}�_��/p��ut���;�0������w�^j�sTmП����3NH��~u�����/���=B��'���pD&3ʲ�Y�p8�>���$����d]h�[��$�B�)Mr������O1D���1�ݓ����5�T{�s�j�'��A���&Bt��Io�l�?�����$]� s(Ep�̕f2���e�;�*1eU��9;�;��);؛T���:����h%��N��p>�,�[��-�Ψ�
�mUSh�m��a��˲�q�\����i�Z�p4µ��|�Y�uM�t�B�[\S�.��f��l��rp:�wL��+-#G��ƍw��\�:R��[�N��RL�c?�ϙL&Xc���0���a�� �1F�d�n�dd:EH��*�.����
F�Tg���
�nS���E��U�ϲ��I,<��ϊ�>�n,��i�reQ��nJ�O"�Hѵ*�Z)Q�)%����m�D+����� �l(��/�lowm�T��R��#��4-��<T���G�s����H������r�艶����ܺu+�����.�h4b�X��ortt��t�ݲ�\g4��65u�U�MBZ����p�xDRH~Bg��x	3
)3��<�/^����}���>��Ga8����
]"���F����j!W���[�-^8�5T�Exn��`~�R��ԝ���,Z�"˪Z�Pt�h\�XC3�ɋ��	�޹+)���8�� (��hȥG��s�δ����7�� �s���������w�e2������>Zg�yA�6�C���6��60�w�ܼg��8���4m�����dk����.Iih�'���a�R0;�����byJ�d%�&��l�����HA�����ڡ�t�q��`#^^�*��>=��Y?Iu6�B"�@�u�$�� MJ	��3ܿG���*�ia�`H���0&;�Kp�P��2M]�N�c���;�B�65�Ǉ��޾�N�a<��x��>`����cq||]�Q(���ƶwթMR>Z�ƚ�+�^'V���z�nJ伧�0�6�K����}rCbl���=��K|!dG�J���m��1wM|�;N<M�00�p����9����ʻ��	�f��$�TPE�x�"7n�����q�v�,�����B ]r�)��h��^xۙO�}n���Y����7����*�������.7o�d�&v�V&J1_.�Hz֯��4Q�[�y�����0��4�y��T�eY1����� Ͻ�y^z�%��	;���O��@)&Y��Iȡ�$�+t-V�����`Z|ݰ����׸�}�&�T�tƢ��*ô�y�`���5�U1r�Ag�L)�A 	%;<j�TQ}C��S��L��F2��O==�C�0��e��˗��e�}�-^�e��v����匧=�P�:��52�}  �4�tk�a��k�	7�=v��"]h�+� ]d�C�"XY/s�X.�� *�BB�il�vL뮅���<b��6h7�2�ېP���u����\�8%)����(�t�ᒫ�B+�U�m\��
j��J��%�e���j a�M�J�07Hɫ���&��+I30�UYᜈ����DY�����^W>�ģ+̷:]�y߻�0�}�"���uNH)�fe;:��8�~���:+�xWX�v8�;<�݄���� ��N5��}�[c�����HJ�Uk�$�*	���6��z�dw�u���O��Ȉ��wz���\k�͆u�<�(ːP�����b�e "i�OY����gU5z�K�yc����p���sh}�r�dkk��\F��𞟙Hx�Y����J�ь������1ٽP�h��ƅ
�w��Fk���9~�G���|��_x�������AǊ�i[�U�a��R�#Ɉ�\kq��A���!J��>͇h$�Kk�o-���#�JQ:�+��kƓ!��N�%W���F�
;�rؔ4����k*� �,c��m�'؋�U�rQ���^U��'\�r����~�#��_�̟}��|��/srx���`��t|��$��@cg�|+d������7f<�X�TU�16½�0*dϝ?�d2����>GGG�eٱ��7Fx�Y8�o���D�΅�����ӆgO+�%si1��Z�;�+'F)e�:e:$�=�6�Vz����:	r���A�=jd��R"K�1�},yR!Jz��:Z*��*�V�=�y�ɳ��r���8�?(�&q_�[\���݉�	��{�h%k��9��9
!8>>��������]��5�Ak�`�#���K�"ö�:lRY�4R�<T��`8X�C	�p0�i������U{ڶ����GS�({�
6
������.�\�"8f9.��-o\H$2�RV%B����5�5�U�"j�"s��`�z��uly�,mMc I�^u8���,��w�mB�Ht��7_�;M!�'��f3�&$Z"�P���c�Ҕo���{�qxO�3�d���ǯ	��O�����-�:�>�����_\���{�w�y�w�y)���ܾ}��xNn�v��^�3�$���d���.eYr||�b>Ge�ic%Ǣ���߿}�Tۆ
LVdxk�#n޼IUU�#�ʩ�%�eMk�ɘg�{�G}�^x���|��s�O��,��\)�����Xd�d@� ?e:�\���������cl�h�1˺�Z�����r����`��٭��(3w�r0�(����=�s���@���9��i����� /���֔[� '�3�0%X:)�S�2�2���jq��C���w���oҶ�+��ҕk���G���;��g��?��?���o�i3)=u�Dy�)h�����D�#v�R��⺮�"<�H�Y�����x<�i�^7���b�~oC�"��d�p8 �n�������ɤ���HRw��,�]��4-��g�K�*>o�mI��R
D�}�닻���ݻj���  ^��yZ')�H�����lk�#��\i���a;h��-!�l�#�l4a<�k��%m���9mt�LD����`>у��i۠��d�XK�gXc(K�-Y��&@ڪj2�@z�*�<�0JZ(��qОoLP���%ZCU%��� ״��\���kc�/������,�LS�KyrrY�Cs��9�Q�%�}��p�u�^��;�݉U�*����-�;:U����5��� $z�Hb�rt[���iLk�޿���P�^���R��FMI�1������q���]ZtEQ0?9�=.^������[�o���`4�X.:��N�lV���x�횒\�n�8�����>����x�"/��"m���o0����P9u�gm'�>�:���(�jڦ�{{d��u/�o2�H����X�k=G�Iwl������6L&�\~�1�z�i^|�E>��0�ͨ�p.�,䃠��Z��>��1A˽"�E� �mY1?YЖKn߸�훷���;̏NB5�X|k0�����o�\,QZ���@�4ت�wn2�C2b�ih�%��%m��?�K0�L���	�J�B������0ؚ�s���:׈<`�������Z0��g!.h��e�0���&���e �e������~�i>�S?�_��_�?�#�����cgw��rLwR"���8ܣ�=I>w�e,K��9�	J�{��\#ʆ{[E���t�|>��耛7o�%σIr����Nw�&��M�\4�0�RhT0ꚶmqn%3�惎_ $�ڞ�vH�S�I�bEj\u��˩-���*?�q�
�9�)p�}^�Z�T�oN9�W�����|y}<��q�o�^~f<Lx��x��52U�L�\��f�YڷQ8�ɝ�iH�Z�}��
���$�nhዮ:7�RQ.���x�����ol7��y��	v�`q�^��V$��5A�!Bw����Y2c��Kp�M�J��p��lԊLp�o����]$ޢ�@^���,˒[�na�AF�g���`�D���I�8k���~��%�y��7x�������y����.���ZdF��.������CZv��B���5�rɲ,JѻwD/�b�5AGd4�h=�ih8����5�C��$Ͻ�>{�I^��G@Vx��A�T9&Z�ʈ��E�@(�8�Be�J0�{RR��9��ݼMyx���[������۶dRSd9���b0��s裊�ʐg���TUU�h�bD�¢G�^���Z�)k�D �i������̏��}s|7�@9�x�䜿r���t�
��㴆L1�3
��\b��U�e�b4Kt����`(���jQb[������'f���y���O>��|��ȥ+�X[u�3���dtztH�]�гB;�>���Ҫ��Z.YV�de��A�G�,[�W�cUU�E�۩z�'���I�X��&���E�睆����F�ogWj��<`��i���C]�87��J)�P2˲��ٯ�{�\���5֢�j7#-�V��׹�h�R�8�x���E�g�\b���4ְ̭����������qy���~��	�uݒe:�N��io��.''s��w��dZ�u�Vz-�	8�Ӊ͊a�{�O�T]�7�z���Y�EVh��?sr��d��h{�h�vEx�.^�9[����	��6G��(ͦz�ܢ(:�@�$;V���L�*���"�֒$o�e�`8�駟�_��ɛo�ɹ��n oM�w����U�UM��~R�������4��u��.\��������گ��=��ѹ%����m��+��ƣ1�r���>{��q]�-݇ə�N���	��������#�=�?����#?��L���/�,��8m�M�RYΰ(���������*A����^������W��λ�e�!�G��t��J�|���BHT_ ǲ���/�Q N5Ɛ
�a�ئ�-��bAkM!��0&�6,P�dk:�6���4�Ҝ�i7�|�b8 Ȇ#.]{���\z���ϱ=,0�wP(��:<A8�*�\��ծM�Jfg)��y�k�>�3�<�'����_����U��@�}/��M�Y���yH:U �*/1΢�m��X�������=�锫׮q|pȭ[���t��S�Ut̼��;��u���]VR�9ؘ�Ⲉ�^U��=i�8Y l�"̎�p���N���b:�`�Mo����s&sb�s��oA?Xw�OS��n564�f82��i�X�߽��ۍ�~��0�}�"&!ッ#����2������#`x)��V5�y���S�!:	,�� {:=�MHp��.BIL�`��t�s��=�p#�P��PUeH�⠓D��Jx�`X �d�5�,+t&A(�Ⱥ�8�q�n���źu�VG�p�k�ϒZ�a8�L�P(�K�Ω떃t�#v�x��<;U������ݟ!��Ͷ��ۧi����>������������.�D�x�yo��T1�Ŭ-&6��Y���Ř B�Md������h���!:�TM�p8"�r
���O������믽BUUL�&��D�!EA�Gg:V�\�,�aA!�
�^K9�|G""���$:�h����Ƅ����l�\�t����x�#?ĕ�%9�����]�g�,�
%�V6 �ˊ��y��q���d�c��7�ce��@���k�
�*�uC>a%�u�h4�5�G����eTZ�)[�1 ��炶�	���\�\.)㹙N�t ��e�����8�Q�B6��Zv��|�B�W�>x�7����^��S�?��˗�p�2�քc�Ҩ�F:�2����� ��:,x\�0�j��\y�Iy�	�>�8���?�_���r��`L''' oR��ˏU`!Y��2������H�#��a]8Z��	ml-eϬC�`�QUU�a����E>D�rYŪ�
Rv������E�?_����\��(��$ ��}X_[�X.kvww����uJ28<:
ЛM%�S;��)�2t���65���LN���TPE8�Hm��4�q-,,�'�z�:T~m�bۖ"�0:�)�ΉS$����ں2,�Op�!��L�G�S�Fx��72��r��L,��n*��q�����В��c��Q�{�.߮�"(�TUEYUlmoq||L��\�p�u]����Xz���E���ލ�	�B��珎���ڊ�)2�ɓ�����vK����}{������$B=|��N-Ʈ��32���Ί�i1y���<�D�^j��k��1t��1_)��@���m�ߚ���gT��A�e+�R�{�3m��599���D)͏������K_�y�?�D(;�ZJ!��A%BD��>LD�5����Nv�iZ��r��9��!�^x�y�ߺ�+���R��}���c�`P"��Z��rvVU$�I�V���������&�pmZGU6Tu�����T�g{��}��y��'�no1��EF[���
>Tz�� @����7np��ܼ��[���d������@e̦#T\,�e&��` z���Pbȵ��b4�1��x��.^@D�@����6GC�u�)�,;2���rYv]�4���,)�'���_,iM���>
A63�NY�1��6���#��cqc�/�9_8w�[�s��'г[;[����P���L20�SƪW>��,8.���nx�g��>�s�� ��������U�t:E*X,��Z���`�g�d������g��宅o�B�Z�.�t���b�k:�u)��D����o2�53�L��3�/X,�sbmoqzv���Ԉ�^��*dXp"VI)�a]ľ��s!}��	!�8���{�6�=�x�κ�ʐӑ����,,�1-֚���dXl�Dj�Xok�+���,8D.� dYv������o��0���0�}��;�����×Rb;�/�h�G,��6�����>��X��Au�+G+X��\�5��βd�H���w�}I_�G楟�i���i�g�|��]�{��HD0%5ZiF�1˺�H.I� ���M�Cl�����ƹ��]�v���˿��^ekk�A^���:���f�	:��0�Y4)��K��(�%y���O�����3n��#y�'�x�"_�җ���>����G4e�%A�?E����9�_���GbZ�L7�&�3mmX�5��O�����O��y�G}�i��b�ց�]d9�(��1��+�'�z1���9�;`��-����h�kZH�Be�7P\*�����s�v�\d��."��E�x{���m�G�M�P����QC���roȤ��t��(���p�h��8c��`,#J �ii�W���}�&�GG�_}�VHL�P[6�^eY���`9?�d~L����՟�)W�z��������Sh�#%4Db�Su�e'��e]2����_���_�<���~�/��,����n�6L[SLgE�bQƎӠ��:M�����N-�$�v��@������d�1��!���R�L��,�HZR������X�h�-
�����4-�qP'xϬ؍HcG�N?g�9��Q�lk�hN�:�~�?<k��l����CD���A�{��:����6M�1��v�#G�b��PY�i����c�wf4MòlR4{뭷�R�����6��{+^�/�Y��䖈�ܬ�n2�S��?�]r��(y��Ƞ?� u?Ѷ�ܚvmp�S"��q2r6
̯��M�� �%p_��^Q�5E�������$��q]1;̈́7	��w����������)��4���Zu������=\�M�g-B$�d�d2��䄲��v�/��eZ�{YF�+�^����6�ј7^{-T\T c�U���`��Ø�y�^Y�8���	�xZ�p��-\��(/~�ü����~���.�'LF#�ŀ,W��FVeB��[�h��ͷy��_䯾�n�c"�gk:���;�,�%���l��p��U�ww�|�*���.\`�=���l<b^.(����x�
�@�@Kj$y&��M�ഢi$�4���+򠼢� ��?9	rMR1��y��3*a�����;�\|�)�j��`��}�����NP�pR�LF#���CL�R-�x���_~�׾�5}��\~�.<v��.1o�aT�xM�P�n�bZ�􊂼��)v���>��=���g���~��^}���J���>Z�x8�(�31��{����L�Nr���
�0'�A��!T�TY���ǰ|W����Vq5Y�7M�o���H|A%��nKH@�#vj��}OYC_��~���,����s(Ҭ��k���mk�ք�r���D��Ӈ�UUP'iۖ�r�b�`wgW�޻��B�?X�����	�ї]�{���q�QW-Y���7ov�]�:�j�L��%B��,fYp�Im�LgkN?��'�BGA�j�����8::B+���AQ�Tu7�J@ņ�Ek�	�,h�JyGr�M�p�A�3(
����ȕ��#�L_�,�TFC�>��4��Y���1��ʭu�R��/F�րL�4U��c��!�D�9�粖�NH�@tk����-��Ŝg�}������/~����|�u]3?>a{:��� :la�]��M�fY�Uul�"���@1����/������G����$�/_&�s&��\�v�,�()���������xD����b�`0t����*w}�~�?�IE]�h��JR75���'���Q~�a��M�x�0�L���� K��iv�#�y�����y��/��ɘ�b�h{J�2���1���lƕ����ի�w����)(FCZ�9h��ۈ�ڔ���dҋ0ȩqx	�AA����ZPm:�j.��bU��l��86��<j6f���8]�
���+|��G������W8�?���w8:8d�S�h��`+���[���ۯ�M�������~��\ޡ���2�a[���5,�sF��������{�s;;<��3���ۼ��W�;��l:%S���1���f��"=~�2�y��J�w�E���Erƒ�@�E��'�=@�64q�*�U4>I1:[k[�q-E[!2>�}b�?��݌�"�&�V����l�R����p~6ȩ�0����g�Z*�;{J3	���F�Gx�YF;k#i1E7n:���<:�� �� թ$ZF'@�
.,� ,N�8��D9Ӷa.��N�9���poD�o�{k�{�ˊ�`@�3r����֨,�U�@��뺛3Ҹ��;�|�������0_��8��x��>`����b�<��(��_�\,�u�Vp�����>`b�V��3J�4}W����-J#���]��4Hwww��tw�=tK�P2t5��1����~�k��:��O��֢6x/��YY�,���(�G�Y�F@�}��/Se�י\h����Y;mo���i	kM1|�_�Ҷ/H29>s¦��QO�����}�'Z­w�w@��n�+�D��0�+,��00|�)��c��}4�܀���[X�P�Ln%�V;?�RP`�pG��L��!?�����V��y�������C�sP4���$�{Z���\V���9�g
�~�������2�ί��A����(��}�o�V���l�x�.\�$�����q�.��2���Vz����팜yq4_�
�g9J�#е��吓؆��j�����y��G���ɣ��	ц B7e�Y>.�X�%3p`�gG4~�z�Heʚޙ�u޳Q���k��`6����?ڂ[������:�sj����v�t^u�J2XAb�ލ��P��/�oCo�ďZ����vd���L�~������g'���$�v�x�z:1)o���[5-@��F^�qf�(��}����+�*�'6=����S���e��?4����p���Fy�X��� �rJ�����zqC���_j�(J@ʃ^z�����a�)Jb�Q������随����	��D�ԢEˠ���v�����KHSk�M��S��FWjjj��.�	��G�u�̓===qq7�|�R�H/Ż�hS��qӋV֤p���(o5���Sl�1�j]>�b�m��T��+p�:.������$�7�c��� �����L&dcrh���5�L�k�%)C�5"�{����gom�;�3�D�t5�����YgH�����ኯ=̄7��S=�|
��#Q��>ɐQ���N�f{�tS�k�E�J����΂;K�d�sT��4k-��u�����;�1�3��	X=�R���������| �)V��ą�Li����Ȕ�^��:{�y<%�w� �hƷ����:�fV6Mq��\�%��N0��vL��{�М��B/�Fn):��X� ^��d��\� �i�+S�C��i�iKa+�)r��˯t�rj_�FH�¼+h�Yt���m��f�VQH�v������V�o����g���i}!ӎcp1�I�[��K��r����e�w��o��-��Xh|�����8
��-��'�#P�8tt<�R������{-��U�������̠�l��[G~�>�e�̃�q�f�����7/��X�F"AH�h�j#��M��4@��d2�\ɧ�`#V��V��I��x���$���"R�c�'8��`��x��N̸1���~�Һ
�(t�L\M?�a�89?0���y/�*�����Qw&-E��='�i׀r��_>Z~�o3DO�b��<���_E�L�y��3j�w���FQOz�Sߍ�W��70]�>z5Z�3x�U��˭NqC�mq��7Ŏ��)����Y*=����0<֍L���������_j�բg���/L�:��TγDG N��ˎ���"��hW�GO��M-y�]����]_M{L�`&av<����*�.�\1\pW�����W�e��w�����}o��ҭ�s��vP�z�$1bο�?+�Wi�9Ϧ=��P&�4�}+p�,�
؋3�c{Y�3^�G���ê�s0��~Û$y����ɽ�<�2�T��7�NY�X�n� A%�6��H�Y6Ւ�S�8�V0_���Ȩk�پ	:�Џ���S=�t�v�GQ4���cN���%΁B�i^��Ly��p��5̜m��8�1C���Ƙ���������e����h�w�H�,�	È,-��"+z�=�E�N2�[y*��k��@���vs:�������`wd+Î�t��c=^�75{��H�%�.G�T��{3v�Vf��
�z� ���*��_�rB���ߖ|J��5ۄr8�ι�m����έĬ��C4J��Ŀ��B�7�6ۦ�������1���s�2�h46���)��^��Si>F�^�5#!�@j)�m��z�p[B"!�#�u�����	o�]�̸筭��7��u��]x�f���_[[U��c��p{���94Ă�
�����8xB�}:�Ƒ]�Xf����s�т.��
�R�G�6L�j��ӭ�������N��T&q�_��8�D�9���V�w�W��Hv���\���ă�>I^�i�܈B�y�	��@��6�?��{
�(rT>wz~?
��W����{����*�ش�x8����H6����������?�����IY�"���ڴ�c���`�8�]�+�������FX;F+r����q����?��� *��v����}¶Ee:���bg�ue�y3��c�����[
�f��<	�X4�̤e�Ό(�C�����C��8P��c��-�*KxS�C�-lWJ-VM�?�˳�8�p�7�*�v��YB̢�@a�bx6f'�v|��t9�>M�(�4--���E�<�'�ה-kwѴ���d7�����V%�$��V�d0���X`�\��NC{HT�� n�4�Jz��v� f�4���V����֑j���Z~ڮ{��^%4�
��
��גRp�x����֓�UM��SF�R�E�q�g��U`O��8'h��4fS�B�|�#G�0�$G���wt�N��XG�]�5�S�^q8M�����$�#$�~�-vz? mǡq�b01��R���n�Z�O�j_2^�c���,�+�m��e*m�&T
��mM
��ab%cF狵+���SPD�q������T�A+����W�V?�8��M���!�Ș\�`L�Q��G�S0Q2G�Ȑ�D��B�+n-�~�Z��
d]6�Y9l$ߩ�K���Ȕgs��_-��	�~c��*lm� ��쩊1����yKA@�>�ᵘ����L�HN��C-G�ɠ4iC�DQ��]w�M�M6�/eR��8D Q���^!�#��-ըgX Z��냉ү
��7��6ʣ/>�KS6Y�M��R����k=�@���R�� f���R�}XE�P�5SDct �0$c9:��D�K�շ<���5Y�um~ik�=%PtZL� Tn�R�R�7W����@>Q�:�)
���F!���49�T!�/Y9�R#��nZ�_�v��Kp.F)w`��Usz���#x�>*#x+��$��?��s�x1k/����3�M ���nd��)zT�nU�vո�%�i��}�oۿ�$Pm���v^���I���Ik����y�N��:�s�Ĳ�[G�V���6�o�/֔�,�-�.:)Q9W���g�Ă�2p������D�/T�ꨈ��7^xu͇WD�`ׇ��P�
���| �	f�xƳ�G��؍D�B�X��=�z�uc'�G�R>m!�CC���z'��^��np|Y��1n�B�AiBfHn�����m����6� �.J2T��2+��W/w��a<uI��s/����u~���è4j�xX�-[��ߪa��|�)������ȱ0G'_��na��XͰAq���kƄ��.2�T�HRtv��E�`�>q}��E!}��ЋpuH
H�:���H���J��2���������C4��3���ja��蚖*ʙ��u�n[��ě��x�>�0_PuȜ������u7�����;=����϶�3��]�R7�]�G�r�����2���Z#�⥼� N���炅��$�+�n2���Kv�}czY��ܖ@�7Ց���iq�t��6Ԅ^<�'��Epw�ri����6ě�\���8E+��r��~�H�|�i�Mv�V��V�s�����b��bĺk��{$����x#�M厎������̲����<��-���5�П�률=�axm�>��|��	��o*�';�
�B��,Ɨ���V�jjM��uÈ[��$���"E���b	�Fb�޲ڬ�O���C=
�"�&��#����2߷.{3P��D.��4.�".8�2�^P��ݧ%MSv���S�`!��-g�������K�aQi�ǵ���s�F�2�u��4��u�(ɋ:�E�ԫq(��*�������°�<����L�`+�~:-�ty������ֆ��F��N�塑�������XPP|��u��Z6��	]Կ���S�x����^��'Bi�ܴf!��Ο�KXa��>�O����:�����'��	��5N�5��J�2WD�_wh���C�ht�H>��
�l�^�kJ��e}�=�󚪕�Ɨ�?L����f�f�����'����I�k��a;0�N���_SX�U:�Em�������Q���<����%��4��l����u����=4#�n��86s���˟)�����w����X�Z��źd?��[aT������?c0��?���h'	�"T��Ή��_4�`n^�0���LXy��e|�Φ�p��UP��MN���5;�sʷ1�kQuϊ���C\�  �]~�ݏ=�~��)�L2���S��FƋ^Iꍃ�A��F��k"��[(�������+m<��g��_/$��
��������zF���=֒����{J�\R���q�4G�]���^Q�������GTq��k�ӌ��hv����z�`�iu��T����{=��;>��L���yő�И{m��VW���D}�ZI�#�w�m�M�DT�w&�p��F�M����vv�u�ޜ��]����a��><. y�D'��&�[뒮"p�@�"S,��o�l�em�;�Mwx��g��Q�����YP��K�.����}v���q�'����L�����8�͆,�vw�g�°�z�y��Q��+D�f٘��sL�q���Pg]�DU�݉x[Զ[� = �ez����݇fNΕy��S�+�����f��߳��������}��zWRhP�I�%{)�65_��U�\z�8�>��霌ˊ��{� � Hc?R�F�)MmݸJcNs�#\!�u��E���ii���W����()��v#]#��v�S
�k\�7���h�;\�}��r�2A��g&Lok�Z��Y��6� GC��t����N8��ЗoC8����u��9v�!O�qr�������C��Zl�6N�L���n��[<�S]8Hu|��)O�<!�Pk�>�B3�B�&Qh�6%����&����l��!J�O�!���K5 ����d�M@
OT��J��%{`����i[C=�MT}�c��v2՘���GR�q�k��L��':����],l�ύ�̈��!���m�aF^r"ʎr�����M�����7�_]�.��K�q���PjkJc%DM���i�o���P;��G6���޳��*ш6�&�n+bI����~��o{���MG��i�|?2���o!XQ���fw��K,�|�
yd򇂈͞	�Bprl�I?�1���L]�����L�O����va��0������=ԕ�iԈ��Y{'���l؞�!�Eu���5e;0���'��eu��9�[ 	�u��
l�K�ڏ4"�Tf��"�9m/*E$� n�Q�w0���ɆW����Q�����`)U)���3#""$s�f����ţ>�*P��]i�u<�<p��n'�@Q�!���*�f�����T"j��8�u�͟��f���$�C�E��\$X���F����6�Kl-�`�B��50K�Q�fv���D;u]�.��B��lu�/����[�A��T.�ٔ#w���v�|��~����\����j�ф�3Je�J)��Y��_t�nPS��y ���ͲT@�ɴ�]1?����;M�O�?�nq���_w�l��idҔ8��cw��u�e4�Iy�
�D[)�1I���VF�3j�'MT~\�Ͷ��vZ^߀f�=?O�ś���1ةi �=��t��nTV�h2�7��1� iT��*@�����ұn�ڰ���6�}��ݳ\�>,��z��5(b�)�M%��(�?��
L�7\�}?�{>�\���z�㙟O�1d�S=�f��HAw�_���*��-��׀�(}��#̃'�S�Fƈ�AJ�yO�!C��]��l{����U����b阎l^���e�:�.��e�������T��o�8���t�]
�H����ǝx���YHN{�-�j��!������������,�&������t��ޕ$Y�M\W)?A'�&�-a⿱r�V�G\aFOO*Ƞ�ӱ�<įj"Y��y>�Ki�ߗh*!���O���f)�\� �l�ϙi��������MA�y��W�i:�)�E}�Uy�S��%��ӫ�|��y��kN�_#�*����*Ն�g5rw5�����+�N�S}ݘ��&ȿ�[��7�с�7i�CC>5#O_���h�p�+�u�
4]*$���dlpu6o�޲J��D4 �Riaȴ��<s� x�y���_��͵�,_�?J���\�.H���'�!]\�I)�B5ZR�f�;th�P���s�[t�i�Ҫ)����Z5`�_�c�2X[wѸ�3��a�j�)�)�a/�������Jp��p��*����4��A�2���`�::n� Ye���-��!�
:��s
��z�	�`��>�!p�ƿ�5����+�Th�2�&��f+ZI��'qE��%޽���2���}�u?����X�k�7��3��C����g��/Rl�0r��A���$�f��yR L4���?����n��,��F��P�٠뮃�ԃ�)߰Zc�(�L	{#:i;i��8�ʭ�O�j�e���u6I&K�Z��ВÁSY��b��2.�����{�\��`Y��.r���z�7�=7#N���Eֹ0r"}Բ�d�mr*�����/F<���"�I�ה��"8��jc>U3_����@5�[��P��&�טoV�#V!�2�'��`�����U� .q�%[[[���k�oe[���+��<>9�"�6��`/��P����,�x�\9tz�hQĜQ�o�@��C9F�M7c�]��YZ�� �Z�9�`{o��Fc-[yjK] �}o4��Y���xqt���k�^t|��|���Cx��4tt��^��/B-tNjŚ�9CZi�*d���L�O}���Q3XY"��:���=t��beE1�aj�>�Qhmt%��w��Ǝ��%]�w�v�煮�''����<���6�9�b��jT8.I��;�l�[ ,M���� �Ky�ߧ�m]��fs1g1H��o�k3����]V���X�v���ec�ޔ��V�J����B��¾��KL�sKR��c�[��M��ը{^e�=ԅ]���d�9M�-s"�ʷ�3I���� w����&.���}J��o1.��
�l��kZ��X��О�D��[�=�t��u��Wݭ�,�O�\�nC��Q�$�u\���j���#w�N�_AV=eu5(	h&Ο�S���d`"9S����g��σ�����n��}"��P\�\�/8�Z7�%�����N ,2�!�N w~���r�������7����)NҊ?����c��O�d�~�H��%2M�Ɍ��Om}ƅ��g$�Usn��U��R�Gy�l���u�f��QPw�-h�Dw�F�k>���z��N�N�P��tGZV%�����p���y���SQ�*c�S��}���"�����,�<
4�.O��'x��E�_���3��k"-�c����J���ٺ��:����A�mul��R��k��k�9���X���S�`?�Hy����>$!�P�Ӌ4��ׄl��� �4I�(
��Äw%"��U���;;�y����
˸e���ܪn���g�Ͼ6h$(	�V�.�:���Gl�Ɔ�S!Ͳ�@��.���=���ǀ6�Z�����\B)��Y(3�`���&4q����6Ev<���B-�	)jw%���r�l�6!/>�f�42����]ˈ+
|]���n��M+�o��e�4}�Z��MŁ96أ-�z=߲q�B����<d��+�8��@��Z��B @�=�]�~4Q�&��)�%�{7�G~N6�P蝹��E���l��.$���đ�~��}�pV�w�����n��E/Yp�m�QN���/!��U2������h��N�Ok��<�V��qe��h:��bȸ����ec_F���7�q������j(g���G] �Q!Bl(>
������?&sgjZ�0��h�*�.C���~d�0�"f?Zj2����	���ߴQ�:2
Ѝ�c��|�W%Q��8����� � ��>?�����J�^*��5����57.��-,@V�1���0����?�
#�dM�G��)a���Pv��q���z`?���w2{e��g鿑|�+���Xmw����p9�.���b\�gqf~~;�97���ďhb*BGi��Xz��Lk��bL���!�aC �w!�b��>N����߆�z&le����ԗJ�q�Z���Y�Y$@�MpK���fQpԻl��^0�~�L�/�~����[v32\���t�u�i�o��^m^F��g�^���(M5e��\��:��<����gg�2��G*3���
���
li��;��O�1���rW�CW���iG��&���A<~S~Z���/j�!!,���<�JA);�t'����T����Y�-nˈ7^z�b��cb��K��J(J5dX{�����H��� �@e4h�Z�%���il���B��^��2^?SYe�m��M�B
��ݬ�
}-���`��������
H�]=>�5&��"�A7ua`��oD��L�^�����x�7�/��
�$��_���s�̓�Pw�UA����'�z�K�+�L@�);I§�Ot�	���/"�ٙ��8��2&��N�^�5�Jn�c�x�,Q`���t�%�wન�;���?]����~�k�e�o.NR�_�׾�*S��;U��?v�v~ߩ,��"��h�9W��0�f�J���y�N�L~w��,��Hӝd�kU�MsO)�����c6)�Р$�º��<\5�$y� n/�h�D�P�,�mry|	zv&�*�7�"8� Q��ڽ���؈�1�P�k����gTs���{IxؕU��W�U�E4IZ�y�J�V.p��}Ò��Z=$v2��j���<���\ݸw��j;q��}�;!��;�$R7b=�I5U��0^Ot��DB�A�`Y;ar˺!��������!�w�ji����?���o���h�O�����_��zot���1��[������1�Z���9��W�ON�4Ze�{��"�Zq�|`����(�y���q��2�'���M���)T#��::����d��D+�N�fE���sY��Zsd
��԰�p�DV���4ycKS�T}L�H��hp!�)�,����۪!�zt�����7�)��#-��ۯ�˚@�Z�lM��MP��ZD~���x:�>g�1�(���.�r��o�&`���� ,ADYB_�48�e2����D=ŝ��� @i-k.��e�˺��j��w�d�����M�ڋ��R�S�_|�U��bh�U��C����j�)r{��V��������k<����-��kOP����9���
�_Jj����ӅT@��D1�ϛ�f@"(��VJ����`��u��0��ǭ����D�]�t8�M[�O:Z�grnru�hZ�����L�-HZ?W��:�b�1ʻ���W4���� ���%�����o���4��ѩ��8�^�U.��r�Ȧ������~'�2]��`�q�{�M��pE�]}-�҂�q2�O����X7��T�Km�x��Ў=siy=��ڼ��An�����0*�z(�<1kR��>r-cW������a�X��oW`͛�M������"�ޠ�>��#4ݻ�F8��t0(|9E{ۚ�`������x�^KeC���W�S��}�H	���o�����~{yy������C��xr��y����.6���{dc���[�һI`��B-p����a_Z���&�m3��B�f���	X���Q��c!9 ,ݣ��@�VvEFy�:}w^�&��7�a�a�""�jq����|��_B@H�
ۉ}d�ZhO7-B��A�$",Q����X����� �<ZB��|Vth��Zyt9��̱%��E������1�V+w�a8h�s�2}y�ӜN����Ծ/ߡR6�6�8��h,J�f�GvTU$Rf�Nֽss���w�WoO�r�i @6�<�N��w�M�k���3��S.���v�����g����9p-��������ͦ�м����	��2h�\����a�E��נ�$�$	$5Jh�_@ȌcP�i�ة��_U��.i���G �~��M 7����;�|3	𳀖�������y�Ko/����W��^���]�wO�S����� ���Y4&de� K\u~�� 桂�����I�Y{!U|��������I{��g���D�x��LoS��'`��x�Cbb30J�VVZj��o�(v6Y�(�ZX��s���Q�.2s��Pw����P�W��bd��@M�J��CD�䞍	Ӯ��(� ��bDGs�|;|�wD���htw�NI3	V�V�;>;��D9ޔ�"��uI�O���rv-��Ă+��=Z�sse_�킈$Ǻ����Τ=�nR�U��ş���a]��k��{Q��<��M"�����f�U�C`	�7�ܢshVhr��=Ӭ�����-餿p�GO5� �!��g��M��������鳈��R�%N(T(4���J�,$r�~�������>���=�4�gF��P��G�����^>z�	���;�_�V��U�BE5'�ՙ�Bf�����N0Tk5!=pa��+t��l�:��j��B����V���Ę��(�?��zeqy���3O�-�MKL0��d-n�g�{�,�ts��D�#7hڹSI��b�������Qg |*�s)���m>�����:��ȫ��Ձ~�s����37�4��	~�(Oc��?��D$��nD����#���Ǆ���y=��u���*�m���g�7c��K���<)Sn���B�ӌ���%�m����7��A64r=��~�	a�Cۛ��xԸwym(L�ڣi)I�5�AN��OM�E�:6u`!Um�m%(-�9>�t�bݬ�c��2���0%@�,L���6��|(��9݌V��B)�h�~#�7������x���-���_6�ڧIO������Kk����A��I�f:T�+A�1u���I]���>�O\�;�N������z���t����'ia�b(�(%����؜����3\;U#�g^[	@�0�F��[�fw8g#s�p�`��O9�bcNL�kh�߸��z�9�DQ����H��ի�=��)���%���m���?�-l��.���6�)\��b'Ŏ�R�d�5䜅�y��r�6�4������.įA{Q��b_�x��7d���gE[ �b3��+ E��?����|u�����CFg�!w?�����A�D|7�(~��C�ك��Y���,M@��C�ꆨ��e|7��7$R�7���)�������7�����`�V��{ɱ���Mh��	aY";��o?*������h��}��0�o��q���RY���+,�V����5��¤�s]Z�>?��|aǵ�F���'����;E�1Z��HH�Vm��9��'ՠ�J�fnr:p���[��C�W�;�O�C4t Ҏzd�:5�^�����Ot��KZ�4C̈y�R%�@��;�b��p�F*�����O�JZqGJ��}U�B:�x�z���ǆVM�L���k��
�G_??aQ�Xա���K���	�
�0����b%��D��0^�M�*���z�𻸵�����aCcT���S�ى9�&'��9&w�絓늩��{�,�i�B�h�����O�Á���YQ$����,�J�2�q�}�Ԉ Ks1gUP"�~�}b~1-b��:-T��lV�#)228�� ?���6RN�E�3��׹T���D|�T'6庩^\�������$�ȵ-ַu��|^�|��y��"�"9Lɉ-ϐ��~?���`�%����cy��,hd�7`�Qg�}7�z�vUB�L�h�J��t�������������[�9dz��W:�YO���M��I�H�u��W G# b���@tf�ɔΑ�46�lh��(^l}8;R�X_ѫ^@8U������������hz�����m��y��Ƒ��_ȽR���n*6����Qs��1�֘Q�����@�8�IO�7N��L�^�u��VS�b���q�ؑ��U�淰�u�/���ҏoٺU��޲V��:�� 7��������Wc�;qJ��Y����v�3Dl�������]G�C-�O*�S�6�"��za{n|j9��e�������`)�n�����3!�lLy�JW��&�½���Ib�P_�R�� ��d��{�5���~^��,�Rkf�9�r�YHi�|�(A!�$[��M12���t�5<N�ƹ���8A$�	�r�����>���&:��o��<&s�Of�7����_!=_,Ňwc���<ߴ�.�
�9���se��JH���L�#D��^d|���gɭ�qi�i7�d�1]<��T/Lp��FF"��&��*�����V.�j��i�c;ѣt��;�����|���q>"Ի��EYv�σ�����ҙ�i�!V�xRg�h(�o	�Lˊ�7�&Ԃ+��d�7��YHL}���+�M"T�ӂ����
�SP��_��tFļiZ+ٳh�'���c6������8G)��y��w�w��Pv-��R��.;��/���a���>�K
�/1&d�R�Fm�H�
��YOE�u�q��q��Š�H��)q1*O��d� �3|%T�Pi`��* ��(.W�����?d��a���w"���B4}��)��R�!àrƐ�^cT�yN�H���)��gu�W�afC`�#��]܊h�sZ��`EM�ŭ���a���-lh���rH�C�a�ؐsV��]�?�ĖZ���VV��BW��"�sx��ԅ%�^���4J�3��l��7�M���&[4����ӿ��n�%X��~��|M���S�4Y�뺆1Ј	0��x�i58��ym	}u�f�e�i�s����8|�:�O�~��&i�nA0h�7e���4.�-g�Y{� �6D($�z�#�$3[r� ��.�@D,�Z��v�+@4�q[���Ȩ77���ې�.B��ņ�^_��{i�t�i�5��D� iS�-��a���1�ќួɌ ���gF�{��U{b/�p	z-4`���P��M�������!ɟ>zۣ��lH	b�WF�-*��A
vb�i}'4|��6���%��M8����}��;�� ���'`p$��}F�]DLs[v�U�������F��w�[�2�8,�PWZ�шϻPK�G^�X!f�'O��ɸ=��b��]
oݨ��i M!x��&��˷1@2�y�#f����`W 	-:oe�M0\S��"��sM��|@	bu����I���%�3�,�8+n�9������d�ZŎ�Cx=�TO]\��J��|3楚Y�G
�Ԫ��*F��5��2��r�;L�m�`�L�>����d�KS|�?������V�#���,���"�ځ]�R����ֲ�QB��7�ɣ��Cb�)�`���(�(l}�W?ͱOr�|A��v��ţ���f�(�ˠeЩ2/i�%��ѱѱq7i�����I�P�s&\H�~2�s=9�xXё�W��%j�l��U3�a�Y��6r�ƾ�3���W�SË́>05��,jD��G�籤W����n��'��5Q�e6��h����0��6���`�-�YܸØ��K�::��� .��ۈ���]��=��H^�u�|��z���nw�_��|�8o���]��Ʃ��EI|�M���(��0��Y��9u;&���=�<|�~�p<<m{���>Z�mg����	7l�T�;�+
;�jˡ��˙z�k����V�w��)q=褵o�U�3��H=���Z��0�TdNWV�����{�M�r���K#MFK�Z�D��q��d�hÆD����e0����`o�,$��0컳M�7�w`k��t4��ȕ��x�P�q^؆����'S11�y��4{F�����V3gx���`C1���4���z�R`�͂N`/eE�[�|��m��j����sV�Y���oCZ��1*����ǒ��%4K6��X~���/�O�wk^X�����F��/�Q9�����߆�uk4i�J�hs���Σ4�����HY�nB �O���
Z���f��0GJ�C���
�!����SoQS�&V�gq �s�oWL#76��:��B�t��Rʻ��>l�$��5nW2�5K([Uߜ`�Om�_�R���ە6�����_�ŕ��A,�	WC��wKI��H\�����A{��@��K)3��[y��)4���P�$�b���*�Ĉ��e͘��㋂HW��� �63h%�A��5+�4�{�D7ӡuUEU���%2��O�*�y������L�ù�֞����Qű���L5���H��򜎪����#���_l��������]3M�ޱ����R>�
�^ �a�I:����, ?����5��b���bm�L�305���K��HW/�M�/�����2	�ݚ���m]�_���}Tl�/(tZ5YjI�ɫ;���-�!z̆&�d̻�Ha䇜�O$��4���w��(��D3�����d�A�[3*���_zƞ���&DY��VC'�+�ϸ�̐~�Ԫk�U䡅
��uN�n���2v��Ox0t'��m�_ˊ�����\a99��U�F�;JݬL+Yk���������z���Y��Q�|ȵs[��s��I\q�]���IMN���E/��?Ė�+�9F��z�!��s�ԍ먪.H��[�%����77>����=�`�0r�E7�W��3F�Lz���$Љ���E���s��R�����plV����_]nu�V	1�@ �-۾�AqQLtM�2�߄��m�ܮCշ�O�JJ��JR���N���℆����|�C{��s��|F��Q�?)��^�'�~N405ܟX`�Qd�r��ք\36ַjnH�R��FU�O�/�#�ņT�=YMS���ǤofƔhd�r�LMHx?1���M��ǰ(}�1$�R��^�nT#�sf�ٳYii�U�����Ym�Ve�hg@���2��={�D&c�t]�Y�'��7oll���+�k�Z�ç�AbV��eZD[aKFWK����f_(�Êh@���9M]��#�?k�JC����7��/�*K���m�\U��)d"嬢�G��$����r�H�̆b�e:��?����qh��/��*ߎB���y��&I�M��0_������>����C�4lX�X7r	ծ�t��G������,��R�ؾ��J!��o� v��Ak�PXՂ#1����Ͽ�
q]ǬhrNGZ�9�ٜ.Sͼ�Q�x��O�w�T�{CգP� M1{d���)�D��W,ǖ�.|�7�����qY��`1;a�]泞+Jb��`_�Z����}��@_h��~�q���X�W��#+!��r��Bz1�r "cDmt&b���L��W�D𮖚̆?��#j5=����y���&�<�a-��c�H��`��)�DؕX[@�o���~�������I�alh�h㦌yӊ��vX)�#u��S3)�s������L�Wi�ɓq�uV��9����^���4�L+ۚuG�zȇ��?t�!��׎�)��>�O4�Zs��/!oG���/>�}���S�e�4���JXS{ۯ]i�}��Kv�&Q�d1<aQ��5X�3(�
K��C�Fa6N(P�ٞ�_���Q�C��b���|/M���S:����R��Q�ؿ�*zZ#n��h���VЂ�����碮�z�^��3ز�u���Ю:S���������r�rq�Tg[�����,�U3�d�'�'���s�Ó;���F\��:�Fo��Y��t_*�� $>4smE[Fb۷��p8ٲ����-\�����]}Qj�[��i�!I�Ϟ�蛙�!�)����Q3��T��Jע���p����a����/װd��A�er���&�i� �u�q�3�����_r��fbm����2��,��t�S�����yN�2�R��2Gb�ѣ�K���A�ĸ3�������3������ɓFY?$[4L��:����7���*Z*n�([���� }�ۈBӌĈ����͜u�� T���~-���ŷ��=�����Jؙ��w������ �@"�/<�]�w�������F���S../�-���N��,i���_�ſ�����?�t�]�<gii�F��R>��@�ǣ�T
������D���AD^�*���pY�TH�$��B#e���,�}�*���xL��b��"��:^-n��6��5ɰ��X�������(
�U�CU�ߺ�$EYTZ�Ny]5��hʢ@� )7q�B����cބ־ʬj)��A�vܦZ�H)��x��X/T�ul�:wnS��ZCY֤�M)˝v��-ͫ�x�>1^����*����k��a0�s��Q���^�WI��F~~T�v�{��֛���,	��PW�6!���)�n?�)��+"[�w~��J��q��G�ҽQlg�n��t��Fxs��9:7�Ν;{�g��㪱�����8�Lj!A!䦴�.K\ DUy�C�	"I
�9p� �|�����;h�I�[L�>���geq�l0�Ԛ�p���:Y6��z�qn�b�v�+2�t��n�ūK|���c�*�q�B[M#)���I�w_9Ż��IS���#�J���~����'�F������Wי�N�q�
�����{�$7 r�.�c�2p"hOt��DQ0\�t�*N�K����u�^FŤq�u�T(��ؼ�
Sknp���
��,���(��W�,��o��`H~i�N����?��/�¥�EN��"{zwЙ�Ҝ���n`f���Ď�hԧ�J9w�=^{�%��._�B0 �Ƌ3)%�$;waH����y��'�����_��f���5���>�fY�L�M���&�S���)vu��QD7Lx���{�~fgf�;M��-�,'MS�8&��l��~�7~����&'f�㘵�fff���ŰܲH�1�uԆR)�	�FkJ%	�'Gա�ze��h4h4���z:�?�kh=�JV��`�Tw���^��g �x���־�RC����;M��y��(c���|�#��[,t�}Z%�.��Я�ik�0���Ih���Uޭ������Jg�H�?llMx���,�����i�����b��W���>Y�]�~)�x?�0bg�G�Nq[���'e��Z�� d@����''m��]]d�H��鰸�HELLLz���j��V�8�����y���`ٖ%�gf���iOtɜ�b�J���V�u���)N��
�+K�O�pv�
��$���\��h��X�a�m�3ם��b:6���ě�{�(3왚cau��{1�0F	
,Y��ZK'd���w������	��!���H��;+UI�֮��W�[	�'��ʽ���D��
8���ݳ��z��^x����79r��ﾋ��܁��S�/���3L���]ӓX��wȵ��Vwk�����%�^{��������s��E�����ql�:|�V+ebj�v���F���Wy��w�r�+�K�����O������/~�8��yI��4Øl�G��F)A��q�����'~�<���d�B�j�zC��O�����>��L[�8��s��+W�����i���į�����s�s��9�8���2�E	��st���T�.�U��YL~Z�Z�D���n6�LMM����t�&?�1�NҬ1��}�M�eie�Wu?�X��cq���`\Q�Z̩�-�y̲�8����~�0�����	�-�FQ�+�[1�u��F��%�U�-��;Im;�ɎM����ּB��D;S@6�=�}u�zG���FH���м��d׮y.\��1v[u	��5H��o�˵�����7��>��,� ǎDNi��%C>KCQ�8�x��)��$��Xi4R��7^{�(�����-E���������\�1�-�b�$�x��/053G�5i�M�iSn��݅\�x���g��3�w'��v�/�֯�M��,gCr�N�b0�)�W9s�-f����#L��������r~�*.R�V�=f1��2��w�9/�v�W��LI3�҈S�0�˫���7-��թ���@b!(A�YBCI�K+L6LL�r����k����o�<ǣ��$�3��\�s��yv؇��B#����g�?��f�3˷���<��?�,i��>�y>���25=E�X뫚N���-� �2��>����|�u��������3'_���;�#�6u2ІޠO�$��&��dh`��>��ۿ��������ޙ�����]^����<��/�;���4E��0���եE�IJ�B����{�O������2�W�\b��]H))����=7U�Z�P
��zh�.%:�Lx˲�V�J�	V���1�)����[�?��VRmY��Dks��}ͅvb>±����(x�ۃ�,�� s�������[(����D�����Y�4�Ơ�B(Y��|Ejg�+�O��0F;CV��;!n�l�^o���I��c�,�� �"��X����`T%��{}��r���ñ�b]I�Fh�uiky.g}��ap�%e`�!��(���!� '%��_��qa�Wp���� ���3�5�J�Ŭ��վ�N�u���Q#"/3�8fnn�3gNy�V!�"�u�J~=4 ��|���IE'ĩ`4��K�m��@��0�R��x�s�8YY]ebj�Rk����������o>�h���Nx[X��G���׆�Wγ��A��d���ޚ�!u�
�K�'�-������ ����^��]w��}<@{j�RB�������jL�4�^|��'O���e���;��O<� �ݳ�F̠Ȉ���ZIV���Ιwh�	ŠG*%�:�&{f��P����ވx�C{f�uS�n�(�������x�ß���^���NQXͰ�Ac�%8�J)RPj������E�{�$W�9EN��3�nqױ�<��8)ط� O|��|�{�������[<��O�v�\}�ib$��׻o-�)�cL`�^��)��P;�y��e�$�),�AYf<��o���%__�����䓟gjr�,�6�	TJ��#i6H��QD��&�3���޽��G��ȣ���~�?���o���_��z�)�s�
&��Y]]! �	IGl�68��]��(?��Y_[#%@f�7�y�c�����{�X�`X_]�*��V��`���?�#�<�׾��hm�������j4*���O���n��J�5/���yٹ� P �����EShC�&��ͳ��D��Q%�J��7���R�ؑx��D�kK)�c����{?�<�Q��pCO�����e;]�E���ז�h���֚bw��T���I�'�z��G�~�TD�t�]V�WQ2�|�e3�x��K�|4V��T�m[� ��9GMF�Y�-qѷ�ژ�6'e�FJ]�QR��������G)~q�}?'ᱝf�$`���^�{�ة���A��y�ni�����u���UOxk����	?(���SS���q�5�ϫ:��qL�3z\�+�v�̋�W�<���Ѩ�0C�$�ٳ�����KKK��C����e��4H~������h���η��/Ƅ��^0�059�]�ރ��t���-�ъ�̪��w����_�F��{t�'�ۿ�;~�t��	Eed��V����u�QF+i��i<����=�`q�����Ƒ� g,����n�\q�O}���N�Q$(#��CD�V�5�F�iF	v���+�������S�+k��dR�+������?�#^y�rk�}���CK� /3�i=���q����~2�K�<.����_\",Y>�g�������P*���/�җ�D�ӡ��dE� ��0�֑��ͱ����"q�h49z�(_|������A
���=�7_�8GG�Q�P��Z����O�����ȭCZ����x�{ϱqe��f���e@���b�'-����O|�3LM�������t���m�f�$� �����(%+RW%�(%S݉�}�!�D�k�ɟD����ɉ	`��Z-�c٪4Q�m��������g��܎mQ�j��m���?o*2�;�Ԟ�7�������k*ņ:�iE��uB�������WOB�g�n�+��k%�6&�лGI��Rz�!�<�p�6���B�lu�3���R꒍�&&&hw:���۴Z-��x?��>�^�^��p8$eF��{�z�G=�[�к�К=��q��4Z-�9m���)BZ*B��|�ϐ�X �0�7�=�(I��0���	e�Y�m�#�_]'��EE����r�=.�x�����-l�HJ�33GV��P2ۈ��� ��g�XSZ	�!:��a�oEȃP�����K�����k��������`��h!Y���޹<���\YX"�c<����k=VW7�����6ѹ�Y����U�_�k���M�/m����:�����_�$����O~�@H��>{v��%����ki�	icLA���6���,-1��I���|����ߦ�%������8�-a���R��#]��F|��_��st$!P̈́3�Ǚo"F���I"����*�oF�lw9p� �=�8�m��h��[Ц±��u��k|��Hm�9���Z�q�?��B"��Q�1?�k,[�����_Kn�Z�-6M/�/n�	\܎�~�Nxo��ok-���7c� ǳ�Պ�»�M�A1Vj��=����m�~���r�=��J9����o!%*��:1���:)6;�bb)�&�F#�76��������KI�dw�+7�qL��cyuuܮG^�-/���)���V��X���� ��$A�1���M�"�M-8���\8��cP��}�c�}��p%��`�5���ɮ�B��s��H�X�0ƍ
�q4e�D�bW�����y��o�~�2sa���I�&�PKQDq�V��bĽ�=ª,i�C�.
0tm�c��f���:��;�ʂǍ6ӔF�$	��K�ľ}�h�[D�7:8��,./ӝ���ѣX��^�*���<2JR���[�������௷�ɮs��J�pL��t���ַX[[���ʁ��ɲ��D�N�EQf$Q��#G�/CF����2/H$�(��$I��9B059œO>ɯ�گ���Ο��r��E�l�����/��ゅ�_�D]>��_a�J��`E����^����rM��v�N�HSFE�:N�)���F{b�F��Zo�(�>�~�޹�չ4�b*EY����R�X�8ڭ.Q�T��� ���ݵ��e�&���jX��g��K�;~��*�e%o���F�����2��g��[(���6(��LQ�v�a<���s� [K9��:�����ߛ[�^oZ����_z��:1��n�u�o픱��~M���U�VHQaYkS1��sq���;N܋���Jm�w�����,c8����J`���դi+G6�6ە�Z�0d�ehc����;9�(��)�A�d���zg-�hD�ߧ,�m0�Mu�6�c�vV�oZ;�(a��(�fjr�{ｗKW�b�&�"�(I��QY0�}򣔤�s�QF�瘢��J�3���F,�(B��9�"'i5��c�s��%J�_߀Bè�CL�ο��I�l�J�NO����Y�6�1q�	�DEh))%��!Lbo�()��tHTH��0!�a/罗��[����_|�ṫ̩�D��L�  ���و9x�|�_b��#�&�p��"V��3�etT�L�I'aT2X^ccy������ǞC�Ѥ�h����F��G�9q@!,��b-�R���e�li�ɩ[��&J����Djl�[-����X;w8��K/q��9��^�9¥��t��^�,/\ř��N�����
g4�hI���K��_�/��<R@��ϰ����o���}��/��O��SO��/���(��$�C�2'�F�&W�=�y������]�B2�"�s��>���6����q����KdE��[-~�o�'�!�ѐ �I\��^��7�p�D9e6����7G�JoV!i�djr�@��$�J� ��ݕ��t~sN�7{{����%�B��!q�1y�#����u+��f%5Y�{]�o ]��\<߯0"E��n(+M]��޴�-��"˲m�6ژ�H�fG�v��틼��X��x-�Z�>���<~����,-I�����ܦ9}���ռŢ,� t�1+Ce��&�*��I�sv�末��{�&�w+���Tj��W����L�Գ1��9W��oDle���js��oW<����$�!�u!^CR��8�ug�NN011ś'�buc�<�9x�q�Ri�259I��cccó�{}�6X����u�4VېU��{��+��f���>��&1�=���ɰE�a"L8���X8}��F�r~r{��{g�\l�)��h�)�B �
B��.nQ��Q,���@)�����	�
�r��9�λ�z�$������Q�LNuit�\Y[�@��y���F�����yBcD�4��b}���8�{?��%.�x���h�Wj�����2:/��"� S�(<ɑ8`r�<�{va��h�Msf��bD��TN�&1b�^�����-�^D��٨I�i+�¹��e���<��c����;����35=�s�O?���ۿE�e��������W������'>I���ɟ�	���7+�
��?�����o �W�����ӧ���$I�G��?���/<��W��?ν�����Ű���ദdA@��2�ٯ|�w�}��^�B�tdĕ��e��a��gi���,��� �0�b�'�I)x��Op������U��{9�I�N�Od��;�{��/\���H)pΓ������i�\�3N6�u�a>�c)�h�>�V�������;ckb��/V��'���E�<՝��H�~������+��Xh�?EYP���ap�-���EԕܝQO�5v��F���گ������56q���L�ZSjM������,..2� ��m-��
�k���+����6�^���z1�&�O?�i:��۝d4�ƕ%�Xqc4Q�����<�s�]�YVi(_��֒Mwb����)(�%�|�;���IϞ��˯K��'"��.��y�uS���+���*�1��cx�������I�-r�]欵ج`2n�M�889ǡ�9V�_�[�W|������9��	��]f"Hh��\�K���8�� �� ,2ӈA�\�C�N��>���w��Ga����?��k'�� �����X�0#r��,�i̞cG�}��Ӝ�����Ӑ2��9�Z��BWVX�جX�i��p��E�}���C>�ħ��������~�S��W�"	��?�?x핗9�֛�./!��O��?�gCq��NRꜯ|��|�_��9��:��{�ū�x��O��ݿ����N����_��W�󜧟~��`H�T��UR�h�ȱ�X\�_~�����qD����7�b��%�Ih08T✥,K�4���<aSlYH�MC\]mݾ��Ì�
2�繗�3z�8�6;b����ș��'!C��Vd���Q�Co��������)�x�qt���/*	�����s|.�r��nll�]�n�G#n'��X��FW����T'�u���Z����f`��ܬ�ڶ�Ԗ���f��bp?2~�$�3�[�-���Fǰ�J�&�y���Hz'B�X$N���i�r��de��K���B��D��h�����KQlwg�VoK�kB�Tj:cEwb�;�����O�&ۓDH��uDV���/Ql��iu�TH#m���?I(V��td���x�(��J�%�st�����ĮY�\BA2�(��W7P#���S"&��8��w�ޟ�5����"��H�Ϲcf��z�O�!0��� y����>Dmd�~N8,i����y�{?���!��λ9r�f0b��"�x�n�����t���ݻ�����ￛx��	�kb��^+I��>��Z�z�&��k:�{��N�dzj�￟$����brr�P*��O��۷��^}���)��~�\����g���c!����������9r�{���S��sss|���/�̱c�8v���q��^}�UN�8A�t:F��z�$�� �N�Ig'�w�����7�4�,������QACE����5�(P� �(�����|�vw�~��)��4ԧj'���Z���c(˲��n�w�s �@������wD��I�R^����n��*@�k�_y����4*��x�a?���{R��R*��
�`0����D��v�l�6������E�!EoH^LTD�<�}�$�Z{<�s�0q�܎	+��R�۰Lu�:XN
��NDXJc���+䭟��խs�D��@�����n�Ǟ*%�I}���ēխ9'�Q���'m��l���`�"#C�|���� �c8�QV�k���&\AA�5�f��z���uN�uʳ���(�^�����Nc���j6S���k4A����[��8�����P��<�8y���p���`b���8 �󜥅Ez�u�Rd�,c0裔B)Eǔ���J((I���_���4i��_"M�%��M̲vy��S���^�s�N1Q�v���|�K_ĥ	.�P��'�J;�0'��N+
���F�!D1�w���yw�2��*݉���i��� �)Ѕ!r�l0��RM�+�\Y�+��C�~f����.yn���j^x�EN���`��KR#�R���O����;�q��f�&�������c��E�DA���� 0��Ă2t�=v����5���5V6����%���h���Q6"�R� �����EQ093M��Q���\���=W���>��n�?��>����y�1lQ2�)F�����8fzz���!��^|����Jr,�����硇`nn����5�z�O?�4���wx���ԧ>ů�����?�w��NV��ǎ3��p�=w����,-/��cX�$
+6	�B譮�I">���o����;Z�N�h���췙ؿ�(�G^$e�� v�������������-���w?Ε+�h5����(�CD����.g=I4�"���cC�@IB�;eY�!a�k�n��=���la����m��v�\���EYa��/�l6XYY��l0<�XQ�ý��
���DYim�j\W��<��6v�����/�hu;��Fu��}k'1���\�^iB
����GQP��J�0���Z�h�2�e�B�t�F#�D[K�&�պPrVYk?�yN��F�꼄A��~!��帝��B�U������m;clk]�y���Y��k0cR
�t|���<���ü�曞,��AXM��?[k�֡*l`-h�A�F'|uʻ�I���$f��eA�;Q��-�Vm4YY�gC��>�p�p4b8�#����k�M�h4"
���
c֗V���?��̼g�;M'Pj&��Ԕ�}μ�6Q%A�����'��
���|#S�S�D��A�'i*I�mh'!���c�9��W�.J�ܮy��w�~��d�K#n2�ɲ�D	f��B	����+���Y�q�{�s�a�hN��&�]<�{���C���"\]a��ʙ�>�8a��I�3� ����c�g����KM#�I�-�{�@M�P���v��X!����>�3*/��("�M�p4dui�0��9I#�	�i�K~��;#eXm�x�<I����qH��Q���~�~���y&'&x��gY[[c{�������K|����ʕ�<����o�����;.\����������O}���$��Ι3��o<t� 8��YF��v�F�K؍�C#<�E�S�Qt�gy�p��1�d��{o����3�Œ�
�(�	���t:���x��G9��[L�Lsy�*�f�(	{(�H�����Nn�t� v������D1��%�,�ϧ(�0�D����2�Q���f����T>���>>�ۇ���)���v3�n6��Ik��}5o�����ia4�� %"���v�Ǎ�uu�h���;�+�q���W^!M�aP%�Y�mc\_/ª:�U,�zx��E�ۡ�h��~��!*�T�`0 �q�x0����|�wS���?����~����4�;��$	Zk�8ĕa!�!��K��r�sL�Mt 2���t�~�ͭ[�F:������*��
��,�DM;	�s�0���W^c���`��\��qii�v��m��HF�i�邑.i����;��I��5I���{/�΅+�@���i��^:�W�=ǉ��н��m�bE�5�ѐ��u��*+���.�F��lH��>}��SP��"�\ylr��ghM����(%	E�UA�
�)s�웒Ѡ�=	ai6S��ι��f'�W�mRQ�aV�p�ar����h���{��"MS����LL���̩Soq�]�����#G����w��[o�ɞ={8q������211�������?�h4�ܹs����.a�277Ϟ��6|�s~�N���ӧ�1�2U��j\)�v`����,�<E1,�+�.y����8�}�h����,y��=�yꩯrꭷ�����LNLT�K���0թ�L$�%�X^�cl��w�ڠde�����qҝh��������9b[d?����	XBz�333�2|8 ���ڻ׉R��2˳	w㱶�t<d%��������[(ªe��#�h���pUI����75���#l��Zc����jǷS�1/r��'x��wY\\���F����9��0=�#�/�꒍2������2�{/S���GC/geQ�e#���X�V_(��ݬ��w� � %�(��{�e߾$����(�X_�3��h��:�&���
�>�����p�\
����8��V���/�@����(m��hsף�Rο}���.r��e��3KB@��Y�U%�%r)"$I P�e��g�����f��l�f���SӴJ8-^�!�Nc���XX^�Փo��3../����Ӕ6���c�cQX�J�m2��?5S�lDQf4��c0 e@#m��r��Q�[�HA3I�y�.Jz��k���ٵ:�~�T��~c5s�wc��f�ŗ��%�?���<Y�3==ͱcǐJr��Q��_���ٳgS�S�u�]�yם���[�i�}��N��t������ٳl�<x���)�;O��5����u+ײػ�U�[����$6�;��;z��������8B�~�u��4�$�������R]�QA�H>��'�W��_��	��,�qDiB�1�N���\��*嵩<#���a���-���eccŦ�^=j��	�P�p�y	�rSn+�V��յ-ﻝ�n�=��fb+�#M�[�|;~丝��BQ�7k�D��t��P=UECy�c�ŭށu�a��^�Z[%Ur�����[@YU{^�ͫ\�S찆g8�xB����LAl#Q����l^�j�5��OB]jT�RV��Em�`��8�����n�@l�<����>�k��J���*y��*�qc���k�Tc�CYj��uA����%�
��\���B
�iPQ�W��C��h���N�ף��D*d��Y\\kufو�p����`X���1�:�������Q����g>���&R8'�V2��YE��N�f��U槦)F6
��чI�XlP(*�YN`��^{])�#U�S�FYN��ӓ�A��0cd�И�;��Ͻ�ٓ�pXi(������*y��BVNmB��y���"c�ۢP0��LM�6����D�M��b#/�yɱ�U҉E�s��yr���hc������9�ʰ�m&��,/\%��N#`ii���IlQ����a �I�H���`eu�={�PjM�$�mx&�����U�8�D��W��G eY"�^��s�~�ǟ����n6��!R�7��4�7C�4�MOT��7�E����n���=ǫ��N��$ISVW׹r�*�.\����4�f)���2��<:�+��~��`@QfA@Yf��M6V7���bh5�,#
$F�z6@p�{y�7�F;�Hq��3�u�ݴ�a�4^��R�/�E�ٿ?_��_��7��S���i���n۸��9�a=-�9��^SV)KYf(ZA���vAH��A�T��D�4m������>|s��1�ls�Ѽݑ�n�F�Q�(J���:���++��#��-�z�ӵ�ꨶ�Q��Y����x,�� �7ɩ�w�
+|+&��.Ǆ�ZC�z]ROR��Ե.v�۽]������#�,oi�W�n�6���/�Vg-'N����pHFJ����� �#3Vې7u�R
��LA�a���Ga�g���rea�0���PA�,E1�/ʂ�,��*��x�*P��9q�ɡCG�����U=MSFÌ���-e����`�9�q�C��~v�q����V
x�d*o-�%���j,��}���+L�M0%Yi��9;���y&v�r�����k���Lo�y̭����m B(�6��@�d�MH���A�KG��F!LNM��F�� T�n2C:�Ɔ�h�Cc�����y�w)�e������\8G��1���j���wN���'�da}!�O�a����{����8p��}�˗/������2W�\a�e<��2=7K��&m6荆7�w��@*���h�0��o|k5�Ȉc�,y⎿�(W�G��&�]oHcZk��!�v�(�|�\k�p0`ff�0
�Yu_y�]��FIO��DMà��U�,���H-�T�V05?Á����W�DY��K�u\=��D�UDi�5�'�A0&3ml��G���g�g��)�W6������sWWp]��EH�-A
o/,+���@�ZMF׹6�1�?:�a,�U�mh�ۄa0���y���j�U2��1��v|4�v��_UT�t�f��V�z �JZ�I��6����)%���7XZZ�?�f�Q��
jk�7(k8C��w[��7��xQ��۷�C��(˒$I��$Mp�2�ȲS5����'sk�+lԆ��	��<��c�ZMz�Y�{5
�aʒD5�z�<W�^@9У�Ng����Ow��&V�P�d�m���o	*̰��&�XHgx����M���)��0�?�\X��y�;�g����z�֯,���;桽$��� H��P*�u���B�[��̩��i����*�!�.-͉&�eb�.�S����Z��X���5μ{��kK,��6�����O��(��a}i��|�0�Y8{�4N8z�sssB��r�g��MΟ?Ϟ=�ٽ{��\���9z�a��`yi���nދ׹���ʫ�x��'�H,�T�fi�@V�SZ�1S=I��>Q��ì*����U&''i��h�Y]]%P�a&1a�nuY\\�;��EQ��������%�z�{"�q%��6t��{���h�)�Z� ����aױC��Ķ���*�[��w�=�ݻ��_������חrscl�5#h�R���B�B�1EY(�Ն(��F3;;���W�Y�-�Z?������vL�������ߪ%�ܦ&�]VI�mҝ��3��z�2�m��G/n_�[0�8��������-���IحAZ��sTj͉'���b}}�$I�x�Rek��׫��&���?�'��ܯ��{��!��^�,��msn��Wy�^��_a߿��a�%~�a�$�Y�)J�8&[X#��p�ݳH����!�ﺓc���ҰGJt�(���$�]k։��{Ba)y��2�mp��4�MD#�Z�joH��� ������]w�x�gO���[g�6�R"K�0�J(�m�F���ڻg(�ۯ��K��F�Niv;�n�D�(m2�����5Gw�n��%O�7���.�T2�����Y�$�,
ν��pĠ�����\<�_��_cvn��}���βg�n�s���dـ��U�}���x������LNM�T@>�)�4��6_��������9��Nt����P����U�4���T���^�󜩩)��`mu!%�^���Y�R�E1��^����4eiXZZ�9��G�z�*�
�r�*/���f��2pG4�&eY 	���2��VH�����ǎ0�w��Xgi����
��2yx�~�a�%#�Q�1�2�����8~��_]A�������*/;��b�c��?[����$��zLLL��kiB%��o.�v|-�(�����뽞�ح�"[V[��M)0��牚p�T�����|�PHe^�����*M�6a��Z������a
��S�f�)�q_[��Q����ﮪ�ر�B=���D*9Ƒ�(��txMb�I�����u���
/����Sk���p>9���@ ��:��?��y���d���LMO3���Q�΂0'��@YZ��0��n�qX�|��Z�,��M^�0�Y���F�c���ҕZ�i#%�@`��±���h0D�6%���KE��@l�[*?�X���ڵ�����!��(
IZqJ"z��ڋ/�M;��W ~�ֳ}W2��XR��+�#��1�"+PH���n��;w���0K�\1�laB�@Xt��Xq#�d�j��hE��<̑�a���'�� �t0N�	��5�T̰0����3DE/g��.�:3����$��Y�V°�f�\(���	�ҨG0��B��;�e����qf�
�z묭,3��0F315E��f�X[YƖ���	0�0P���)��k�`uc��p���q쫦������+�[�׭χ���S�S���q��Y�����ͭ��3�sP��h�BIV�VY��hOL���'��0B���G�"JL����(�&N$i�˗�`�#�"ʢ������o�n&;]�I#%�{��2�xk��ȕĦ	gW���ӏr%�a���!'�� 7��hȀ ��j��6��K|�;���'�$IT���:>7�RU[�!�N��4ƖX�q��]a�7q�e�!I#�`eu��Sڂ�=se�T��#�┫�l���5��9�΍Eƛر����&���lC:��5Nb;%�jD�E;�Y87�c>ȤBJ���"X�EA�cr��F�(�@�9`Q�3H��:�M@�ͺ
�d��K*����8�,J�<�s�u�� �#���^W��(�:GE�[�h�l6kr�Y)�?Tܮ��BFј f����bȶV���8o�ֹ1q�9G��q�T��z�Ç��'?��7�x��W)FY��ZVnka0v/{?/�:�ֲq2�H�]����X��@I9�v�ɯ��0<��ѺDX�k�U��u�Mi#e8�ȣ�BkMZ	�+I1�m�8��븢��0����4�mV�CՔ����p]ݕ�K�I�2N�UZ�ƐI3�~�U>�p��i$$̈́յu f:��6��h��?0����p\|�mT�27nc[�
(�	*���}<���L�E�*�>#4��� C�1"1hd�+3T;����ꕫ\�pQ%q�knk}�n�j��o�p�'�mll���¾}�B�իW�e�5��gϲw�^Z��.Y�X��j�+W��n���pcs� |���eN�:��.���q�
�k	T���7O�䥗^��S��3ۃ��'?	���
o��&.\ �c�=ʑ#GHӔ�`H��~{4qua��h��w�MQAH#m@���zlN�k$����"/J�:@��
�}7��\x��;��r�4�t>��� Ϭ����'��w�M>AS
uN[;�&��m6�v������B�E���Z�'�V\��5�t��Tjk�B�`8��l\C|�Em��� �b�m�c�����+�!-[7Ƶk����������F���m��Ơ�b;���}�Vg�FG�g;���ۥ�����`@i�:������S��g��,��.�ϟ'��F�IEt:������=�n������U�ˢ Yf8~�q�
1�B�6������d��ֺ���6Itֺm���)�A�'>����Nw#��VG�$���2�TX����?@�l��>NV�U��׷�n���9��$V��+'�z���M�Yz�Q��XWs��ltbp�^9b~n�C�s��;�F*�T�,T�h��!�E�љ�%�HI����0�̲<ڠp���`�f��<C+ �^�3;v���^z���>��>�1�������Y__G�3�<�p8�ҥ��s�W�^�{���{�㬣;�fmc�����w���ӧY\Y#J<p���9���8o;CII��<�Ѓ��⋼���<��4���8o�FE�ϟ���Y\\���p��IΟ?����9t�0O?�4�7_c�޽�>u����_����Ç�.�s���[E��C����8M�7Q,s΢N��w�sW��m8�ʫ|����F(�bP='�F�����~��17 ��1�Ä�^!�[i��"DTa���u�n��P��r�F#��6�'?���6)�k�Lt�,,,!κ���[J�1)oO�aR�6�5�^9O��V���OV�����$�eT[M׆[
/�Np�;�5A
���ݡ��=�;���5-�^��K?�~��Vr��:3���5gf��t;�wI�+
E+%��E�JI�Bk���E�0B1����('د���.�f|cGH����}#�|�~��'��8GIY?gQu���k˩4��³����x,K"4f�Kn'���}��v�2X���M��q!����H�S�$g?����v���X�+�����6��B��SI��m]�JG��~����;���h��LvH��l�MͦFn�寐8SD� J��"��ϓfw�_wVLnPH�XqC"��<+�ޤx4<��� ���.�[��OI�HN�{X�cr��#�_�A�����@�\6k��Q,���d�G����, ؿ7��Ҕ��+޺�b%�22i����ܽ��dL�^]���B���f%����!>oQ�%?-1Gؖ˶FIF"
����P�2Un/Z���t��^_w��X�<E�x\lf]a��V�`cRb�9k����>��K����y�����Zw?N�â��{Qx��y������s���0��wrtL���:����%����?Ğ����^�2S�����{�ܐ��]<�*���V�����P�.����AǊ��P�4��to�Y��X�ٍ���c�(�r^�6~�����L6�!�u9{[*o*�����L'�l�h��!������w"U������BR�c�$���z4�4\c'Yyk�vWH����a�������RW�Vɬ�ʮ��.9��"���V�s�N]\a)��\^�t��ٕ��PM��cE���B~�.|[�!�x���u)�Su�Gk��T�u,ӄ���;���13 4�F��r�������ORDDD�2�!�D�妚�!3`c�@@$B�&��5f�+�g�lF	�am�Y�k�-�#ݧDV�x��J��*C')zc�Z�4*R�e���~�=�n����ݖ�9[ѳ<�p����j7�j�+�0�Gh�[E(ȃV�`���l6�Đ``?���x��<��μ�,��3�i��ɯ�!���UU��S (����*�?�N.����C��� b�� ������ׯ�����E��re�K�����Cy�ys�Q���{~G���ԫ�5�c7��� ���m̂ӄ֦�ue�ƍ�a�u�+%���z��;�5�GOX�OZ�``.�����a���|��2�}}��5q����a B�����n�������g���c̒��F�d�5u5���"is���H�g-����tSq�������v�L����m>vLN�1�L���v�lH[?}�����^��	��rpp��T�6(���c;uz�A�B�?�YfC����N���5()������D�JʉX 
�C*Y��~J��J�?\7�Չ�h���c0�>x~��,�������G�J�Ɣ�x�V1�*�ޫ���>؅&�ia�(�����\�#�X���e�*  �j"�A�H����.��ݢ�؝~�xF��Y�Z�"���A7�/�j-E 
6�|Ҫ��ZE<���S��ϧch��u�_��a�Hؗ_��_+o�z"hn��^�c��Gޥ-�1�_��D@�D ���j&H鴌��ڐ�F�zgh2;�i�r�Y$�=ւZ�{�"�>9����ވ�g��<����^��^�gCH�y�&3��Hc��%�ܡ2�������Jb(�N��d7�P�i	���- �̖����/�U��Y��}*rL��h�q���%oDs��2,[���<�1{,�p�'%7���cM�"���ESK����!)�PSQG/��IЅ\�tU��;!�<��sM���'e�HF[W�wi���������+g�=��y���B2S1��������njz���y�Ci��؜�@����?g�J1�Ϊ���=����Ӯe����_O���3�O���	Q����ƿ� ^�J�uj�V���VScI��y{2�DQD�)w�ܑ�2���{�l���3ɬr�U+.���t�v��+���󷷇ݍ���e���>�`$�܏G�_&D�.��`��Åݾ=� ���P�ȍ.iJ�l�'_��܅�_�Ѷ��4��RJz�ͯ�>)2�u�k���د/��f/� O�%�6��z�6)�O�\y	�l��^���������<�l�ZScA�H���rO������0�^D1;|b� j٥���\���~��P��e}g��l���t��4=w���Dރ�d㶒lU\�%%��v��;R�j�fcQ�@��wk�~�"�]�<���!� �(�>�~1��ĉ��g7�h�w��>�L@�r���5[1_� ]����s�C��1~z�8�.L��]�o<=9���wbҢF���D%B ƈ)Z�a`�y�,��=�2'.w�>U�hW"���4=^6ѲI�Hݦ^��z���ߡZ��;�w[L�I)�]��8MĒ�q�0�� ��G�������qPz,���ѹ���j
���1oV[;Hd��q�!/��Z�df�)f�}wb2�i������j�|^��d��3n<=@��NQ�E��3	S�����v:�a'��%WX�Am���_违�t�{T�bD⊖֛���|"�s�h��2�T]��z���xG��=�c�^r_(���.���Iw��(NNN:��`7��á�,~�rS�*N���~�;��4�Х)�	�/H�=w;f��ш9�ۦ3<�y.m$��4���$����~Z� T$�}[
C<cZ�f�ᆐ��ةI���X������R5�>+C������u��X'�ƕ�4m�CН��.VƍaH��#�Q�q,�^S;!�/	��J�`k&�e�L���;�\�Ng�Oo�g��P���3)\U�t��PBԢJ�;�I'�j�3Nt�P.M?�QW��/7��<ߓ���+�'�6��T�1ƻJ����.��Wwg�l�^��A���,�b�3}�� �
c�)��!��N����.
�n�.�;:�jYF_k�(��~B�6(@[�40}����߉^�`)X�Ѩ���4Ҟ�������Y�e�u�Xg̛>ޝ�*�r��E0���S�߿�^_������w�eqт��J��:����W|��1SM��_m���wD?|�M�|���I�/*�4�,�C�=��R�)�d@r�Bi[�Y0��_E��cU|�q��f��N�G9JzzN!>������œ��W�U���v����Gυ������E�W׻?+#�Aa]cW[A_��A�cN!WH>�������'Ks�"{^&z�B���Q�I}o���ʈ@jg��Bo�}���s|�����l5N`lN"[{��FF�}��uU��0�Ѣ����6�mH��n�bu��KƎ���H���"U�����`t�]�3���j�h3��-_���P�p���x�1�b�Gnҫ��\�6����ޚ�"���?x�p���?e��_4�g�.�������U�Ҹj���6"�L8��4z�_b���5n��d����-�f��L�Dg(�l�w-=N�34r���Z��#S�{�/WlzSu:�F���э�s���|Qu�[ШZ3ZR�N��M�����
y~_3z���o
���?��I�� ���G\��#�Z+(�5z��y��Fbҵ�ŕ�^��Z)*�r�w��G݇��i�^��.�d�5o� '�������Q_՛��7�c�A��T*��.2���Q���@60�ga��ϕ�7�&8r�R)����>
��ݰ�ֶF��i��x�m�4_�L�.;V��.<�Y3%�¨g���#E�����1d���MGm�mJTXG���	��t��:/(�Z%�l�����L��S��!htS�1��nN��p�A��צ��4?��^'�66~�Sgm�<g=�%��<�@��<��\3k����@n���D%%L��S�Y	$�jt[ݲ?:�|��FL��I�J�J*C��HC�3jNA��`s���a�H��7^M@�o������x�w������=�%}�|0�ό)�'(��qy����S�����D��o�9��Űc�n�Hb� ۓD���/�UU��D�k�
�,`B]ͣ������G��
��+�E���%S홤GmL�@�qs�{�R�#hZ�s�`��}���T(4���X#����d��7��U��'"=��]�������N�6�8���#��DֈC������̗��E���$�-Tq�.�i��a�����VsO�S��\LK%,LwDr�<9sN�3�
��g"�oVK.�#G�P��G���{�xF[@Eb@�BG0dU�pY��H���~f(Ӂy%VI�ʬP��������I.���I���>?bE�r����ϭ���0�U͡&����.�b��_,���8�l�j��|V�Q�m�᧤ꕹ���C#"���f�͒c�}���;��p��m�劁����/CuUE�;G�x	��{8#R̭`���j�&	�������=���r��
D���%K�����7sh�J#�fМ
6��YC���KY\h���-��O�Q1�TqE��+#KO,N�>/1�@Y���9���C������ܸ��n�sL?�\�%��2^��n�wBC�:�9�N[��R�<�`K��u�>�Y�Ϝ4����|��[_����3)�wQ��^l�1e���k�8|k�	�D߰E�9��M�T�Fǡ?�?}#i�Főԇ��<0s�����i{U�G{��7�R��!?������c��g�ICW���o�gS���b���b������;_��U�㢮�U�w3�k�U��E[��:o@AĎ���?��8�C�A:��`cW�t�{�z�;��Yt�Uؙ�,IDO�غt00�<S���:�,���K���RA4`�t��+x#=�B��A����y%*y:��S�ڑ�S*ӎ�Ȍ��R��m6E�5���\�b�n
%c��r��?Ѕ��m3-�[Qn�Z�����D C�j_������4��`L�S��Z��Yp͛�ve��Q65���ʦ%��ػ0���� Ē��)�V�����L���8���ۗp���ӡ�� ���i4��{��qJCt'Y�:C�����J�'_(kAr*�;� C )�/�ou�~ř.���'��4D�%V���R�&խ���1��������*�m@W��N����a���Y�7);�Ǆf���:탧7 �u ey����\�(!�I>�j�	ܯ�/l��vF*�K"Q*GG�:9PF���q�ZBe���|ݞ�-�b��؟���6|k>{M�Ϛ�� D�8c7?R���3��ݿd��S-�sҼ~�ٓrߓ�	����n*�;��{�xy�|s��$s��,7��m�H�ƕ{^T�����;�K��~cmM�V��zB$C)`f��2��2�J%y���Ȓ�m.�ߤ������%�R��Z���cj&`�u�kˆ�:��*L���j��nd����Ԅ��M�
��+��Z����<HS�X������1�H��~(mii	�	�Vh:�e�����F�w�H>h!�8_pؽn�6l#+�O�[Ү=c2Y�k���)����Ρ�v}Lc���}����l7��!�:����f}�~�O.1x��X��On�iRp�u�7����nEl	��j]bꀍ�j��	7�������D�`��^�TF��6���,A��-JD;�YUm�L��0W��a�F�`������aB��Y��Q�p8a��\O3X;�_�KE����*�sıS���u�bbBSa�ؠ�ADB��l'CO8w� "[(���'��M<M�n�ْ)	V��ܦH���6e����4�ty���VֆK+dQˆ
aaLU���?|]�4�L�_J��f�*�gRT*y�eg���_�;n�~�~��wz{��;��𩄖��yC�8��eV񎟗��ئ}P(&22r��������y��NR��E�S�gX�ÃL���7�,�:�g����xo}T��+Y�N��̤�֯����9���2����*��>PF��N�`�^�.�_3'��)�'�˯�36_/������)B����2Nt�~��}��yB�r�+~��y�b�g�?)�(*OJ�mwF+���I*�_XBB��y��&ꨏ1��_����Q�zk��|��jq�Ѣ^��^��.Xk������-��}+�2^Ԑ��.� ;e&��
9�|����*赐/����!��I�/�|��Y�U��' �-��ë�6L;�=�����J�x8.�x�ͮ)C�3�f!ԮEV7�4L������}�J����J�7��G�Tr5CI��_�L��/��S$���faW��,����i*(Zy1ZW}e� (E	�ա*`[�cH����O�7\��fh����[T͸����e�YٚjH�_��n;�z� e�cα��ߥC�/e?5*F8f�iF��٘bQ,��ȍ�����u*��4�������,NV���Iu��)v��q�D�veԆF��m�v�L~P�gͦ��^*��jԮ��C0
�i��29��� ���d>��z�]�0�\@eYj�;��X����.�883�꺫�HK���F�,��6>}����o������L$}�zγ��C+ �1+��Yޜ�}�&e9�e��.�u;^!sC���e,�~m��혨qE�E/O,�t��z@Ċ(��3	$�/�C?d�����2��ZȢ���+s.�w��8� _�У�a(�c`��ը��io�<�%leW�\��忝���U�UHx�#�^1�3`�(鿝6s��_���H��|6��L\���qK�"�5�2#��;پ�f0x�ƋT����.Ҭ�g�]>C�� �!;7���\;��E�ۏ��H��64ڗ����l[N�֘�ײ��K���<�GH�ݽ4P��ԲKK��b[/?|�#S%�����@0\ ^Z4�����.z90wU�mvDK�B�d42���OM-��d��A�҂3�rt�����P4�x��W{B/
�d��J�O�D �7����,q��@�ӣ+U���ʢ�}ЌS�]��0-�*T`a	'�Ռ�"�;6T3v��Uw�-���W���T��d�f`	&(I1Ļٿ�DbP�ޕ��vQ��g��N����,�'G@H�L� I��ae��buT����
ب�K0%D�4�4-��L�@�b�%1VZ��{��[v�cǟW�]��f������}z�I�4��y�����E������XI�A�0&���7�$,�U[4���IΤ$e��E��ׯ���u31w����^���n��.��]􎨈b�mniW�{�5o}�����Јy�Y�~TW��H�)�	�q��=h1�5Uل�y��S��� ��/�k���XZ�L��� _FŖ��qZk�-�����~U�|�j�?��\����I�O��aEk��[x�F6	�޽=�gNC{��<yE��-M^�uu5F��vf0� m
��4XI�^]���;�b����v#�O�Z[�5[y��A9A�V��=��DT�gT�5�u� �����R��k�A��o��Ѥ��0N�ɤV��W�_PW�k�j�L%�	Y�߈�OSf}T�T��\��8���e�gBs�8ܴ����C�P���M� b��D�����/R3o�(�ڬ���9ɺ�����ȤD���+b�,����~��Mɳ�{���Ԙ��%J � ɽ2��2�Y�����]���b"�}|����o�e�n��`��\L�/o�]�+�n�G���@�]�����1i �Z�[C6.u�b
�����|���|�W6US_��O8ĊZU}������u���P(�F*�eͽ���8��(�mJ���h����e�K,� 9pP���*�@��ޖ��e��)� >MN6FP'�$Q�����B���]p����K7�0[2B,ƕ�vVq��vȴ���H�bٲ�-��o����ӷ:ȜMAU���������JFC�E�b���h)��)�¹�wf��ܻ*�����K�D������(P}P����~9��w���fQ|	bA�hJ����CV#��xޛY�C�Z��Q@�E�Qϳ����b��-쥯
��`PU-g	�&�P"_G+���݅�w���ǔʯ)K#��?ޭj�X���Ϣ����	M�E��W	ς�ca�5��� ~¯f_i�J�����,���P@$�ЏG�"�2��q�)� �"�#���g�t��>-ٜC�k^0�E��x'Z(��\K�"����-��u;�6�OL "�9��ͦL��vN��	w��^�!�_�@RD�r�0Ѯ2ţ-�͍\������i���f��M6F��cf��>�B�� �ۧ�7i4�)nc�ٳ%ҍmpl��T0zq�nw��Fl�������V#��t;g�q��~���'�j�����/��5��}Ya����f������Z�d���)U3�!5��4ld*	+�=Zi������_��*sKN�l�Y0�F�f����nb<��5㠣6�ymI/�x*Nʹ����c�n@���T3UI�����`e�x�%�S'�x4�XSw��	!��gN��|&����4����8�,^��H7x�R:3�UeT$0�����̊=Ke+zH��j	�"-~w. ��<�O���fL	�#����#���au'��,�7��Ŭ�&1eNf�EB������n��>���"�`B�����+�VŌ���<E�X2��������7ò�P����
�Z�4ZX�dbS�a�A��BxR�Lȼi�y�%O%���(P�?�\����:v2��*��S�I��.YîW\��"m��K����Ey/륈���ޖ���*�}�*���-f�h��[��V.��䚼���-,�m��F8�yoV|�Џ��Y�����P`xr�X��v��ZD��i~98���Q>(6���b�xgC��`o:k�����o���0�LTh0�s�zz�^^�D��4]wv�1�ڗ�(9#�j������\ܿ��U#�W4��бB���g�)����6;v��w-������$�q�a�Q�'�o�?AC�5�+@��'��u����[c%�ŗ��/ݗ��t2���Ź���qZ���^���i�O����oɢ�EyLHL���
*{��M(y.z�K�-�]]^�֠�JU
~yMwp>JH�͎���$�E��nwOD�U�Jj6@���i�SL��-�m{�6�¡C������~�����@f]9w~l��Oψ��11�;�fVN�!!��H�~�H6�qXA%a��HYEs��#4v�)p��Q��F}P�����_+/ �_�#Q(q}!��Fc�׶$
�y�j�،�n�X��THZ�&�vv��`�X��]_�Yok_��C�u�E!��Za�S�[�6���Ħ�Ke��X��v)f��Z3���<t�*��S*6��n��ȃ}���Ļ��Y�<��!�����1"!E�Z]j�xή����q�~]�~���Ȕ���f�O���?��~�6XЎ����j�PG}�Bp;[(��@.Y@ܽ�	�7F�p3[�/h|�������������}G�`���H��5��bo�f"?�Hy��%����q�z-,�[.q��̈́�������h���g��~B�6����Vua����ȜrF:,Z�- �����zk���:�4-㎏ǲuk�k�p��b8�#Ȧi�>����h��fg��S�@�U4��8�������ƪ�}<o�33� **}#�i�l����p��6���	1�թ���b��]l�Q�RV]�Z6��
HI�b�WT��'��~ɗ5�/Me�2�0���"gp�]bo�K��������}��X`�j!ƍ���ՠ���Քc}�ê�S.u����Y{�̨E5d _��Zy�v?��bBe�e��s��/�d'v��|j���C�#�L��0�PV,���i�c�C_?ڞ8�½i2�8�Ƅ��9c��ZRf!�Oi�О�+µ��Z�K����y�dt�ߔO�_A��������D�F믆����q�)#��z���T�����/�6���?�J�B���(�����:�g�m83���4O�Kv+��bS��瓪�ǂ�z!NZLW(��E��zktȁ𩀎�	��oք�wT�c9�z�{u]�k���j������M�̤b���8L�{�pp@Zb�]˰�9�1�JÜ�F�]F��R���%�d��N��_L�V�!~��ڸ��Ut�������｀��c~m����8�|�Y��d����ܔb�=��N1�$!d
�mm�x�E�c����=� �G����0�#BJ0)-hJ'?�g�
0�T|lHt����+^H�n���Wɸa�����Ѱ��ѭi��WQNA�0z?������wB����>��}v�����\�.�edsK+��`��%�����<�t0��nќ>r���=s�� �g	�:���P�e������+��n��':e�:���"��Z��c�̍�{�؄Z���������j�ko+��m�>|��fs�=#�,q6"������q�WC�X���{$R�ٿ��}O	�9��(�n���ٺ����D׊=�w�)�薵��#��v���> x`}ZEӭ��<I;��Ř\�aw?��⠄R�A�a�}GT�z�PHiNx?+�n�^pw*}�ͽ{�j�9�
��-i�Wd3��o��c��VR��Je�;J+�a�W3;]�y�Cp�ݦ.7:��OQ�ʾn\j%��mP� �JFDV���Ӕ��E��2x�*�v��4�#N(���Sl���48�G75\:��p�@��R�EMnB����n���a���U-K9�FzVS>=�AԀJv[kƐhG�՝��TVn�^���LC�bQ��3Ɂ���k�OB�`�m�~��aHoa������F�M		�*Yg�ڰM�j~�ӈ�ʋ�P�=�!~������m�HR�8�᳐M̽�[!�M�gJ���VW�����}���MBף� ���7�ON��D��J��l8�	E�Gf �ۄ�������A���X��n:�pD��b��[#�q���I���J��0��*��E׌�K�~��e�6T0{rYQ���k��[���:j:�A����诳Gc�[�`"�+V��V)���I��K*��=�q1��j"g5�S��#��'��Mi�D��p� ���*F����bDb�.�<uh���ݛ�J�I�9��w���D��j�]��&�$v��;�r�~��)���c.O�[���_]�����Lډ eU/
:�GJ><���<a���oK�Yb��m2�_N��=�7��6z^�}�>H�(��{=tGQǀ��>�����8�{GHv�#Ы�J��@���*�YF��yXКi��i�CG��#�,��ԉ� j͂�� �
��_�KK�v[u��v��h���	L=W�Ğ�'''��i��i�E��V8�#�4ÿQו�A�Ri��^�A��C_d�}3a��SL����ŊN�-$� w���ce��f�jCt����+�:&�T��7�Ĉ��?��AO�Ù,'�C��x��`����6J�،�ɋ>l�H�ώ�a���|�͛������t�{�g����7�\��`�q�)k�R1[k��5�]��*����v��ő8ℿ�z����d]H��o7�!��F�Rp�1��g
�oF�F�+S�ֲ�E嶼ʘ����hP5(/�6d�i�wYb�Ta}e;�S��'ۼ���U�tLI1d�Miӈl]��_��x-hI2o?)�������ʅG�O!Q��#g����\T�g_�ʕ���q����:w����K�އ�*H*]����܄�ѐT�ʶ�Z�00�����+k�<0�����\�T��˅`nݘ�B���8����J��|\C�ׇ::��_����2��H��`�_䡔s.�x7p�G�lBB��j���P.^�j,e#0�ڢw=-Ŏ�S�X?�,Z{�g��HN鈊,I��P��6���z{�h�a!N���
�3m%�sZ��L�\�u�쁹��:	�u�Eݗ�P
�����)�����5n�m?�۳+!Ƌ����㈁��S�R�./�hѴYg���D
�"��	]��t�FU�2��I���~/U���fHpG���&[��C�x�F�3�t����E����X�O��Q�U=��<�t��Je}��:hrF��V��KV�Ͽ 1+�Ny�,��ə�]�cR�M*��z�'�O�L��V�6cV������9KLW�D�.�m�#%m7�xN�{뵎@у���=��w�+�sU�s�%I=�SP;�WYC�J��(�B^���&(8�>FAo?�4�G�(H��?�u�&	���@���!��@v9C�Ժ�v1C�
T=�5�xl�i�L@C�n���m�u�.���T�N�DU��'.`���\lvn�d���6���V��y�O����~߂���fb��||������kQ�p�#�D�7�)�����!RǼT�ꬍ�|�4�۳�+��&[�ٽs�CP�M	��yĕە�Y�����Y�����-·��7~�@���3�Ϧŗ���k�Fq+# =�����8�L��x��q��r�?3�'|OJB	����8��-5)F�F?sU��>f��s�l;�C�fZ�Ő@Ř�.e�#Q<߽��z�K��̂��:�p�}�E���'^&~>�"�Pz�����_d#���Ҍ7i�����YzF�B�^g�Y(��Z�`�k����v:�y{+��j���Y��1��,�U �Q��Q65��(8{n��_p�4��2ǵ�z�~v!�{�Q�)��C����ho@
�`��+ۤ��e���aP-ʧ����y�a�#�g�ӵ�=�8~�d	�/g��o�-kZ���<N3��^0Jk��3�蝽-��=KC�P�c�#�@�8GnCg��$88]Z�ͳ��F
��גR�o�Q���Έ8�G�nu�~V�RF���Jp���# Ѓu�dl+�N�2N��B�A��˷����;�P ��q��Y�8�!ۍg@xE�@=���^$R�Q!�	㭖m��_�C�,�� ��?���U���mBeF�M��B��ګ���H�*�R��pC��S��|��jf��r�z�?����T�@�k	��%�zkGn��k7O��*�6�	�  ���/'bk�3~�.�/3��$c�&ER�ރu����,��7��ٚ��Ղ�@b��~#M�t	�S+�xF/�Q��X�]�s��`�T�)ƀ]��t�rp��n4�W�J�!��m������ŝr�6F�?���(���ƴ�SR�@z���UF�0����)%�ղ5� �6\B�剭�TRt+/�
���d�<�ڴ�T����7a���2	�3�}p�B����"��~��.�5a�.-C�#��.��E|��Z4�������������?9+�+U�٤��Fy������=�U��A��mz	��g�욍��Sk������_��Cyc�8����C�3e��M�����,͊i���e�w<�o�
Y$��iX[��it�j���?�E�~���g����S�T��}@EE�'ڕ.2��1K�⍝cH�^+k��C���6g����a�NGe�BMw=SfI�#q�;Q,k�3u���+�''�S4A}?8��kd&Xj5G��zU�eM�8h���a���D:�'SbPA"V�ZՎ���&̛���X���3���͕�r����7(�̗�qZSǧ ڟ|8���A�qt(��L!ՇJ�K�;��VMl�DE��w��X�ֶ�)�$%E��]�f��bVJ�ľ���#�|�0��y�,Ao���x��˪j�F�c�.f� �2�z�Oo�$�7bV�G�!�Z� ��%�6���r]j���kk�C�u.���oӡ�ǂr�{4�e��bzCl-�cQ2�-;�A�c}��WX���i?VLI�w��I0z�C�X�,��?袿���д%���a.d���T�#cx�.L�l����H�4��t/����&*��+�fj�t�w��<�p��jV��V;��uv[���_�^��<�qc`�EDD�����T_��	t�Bt!%�[O5�&/��k�gM��4���5Xʁ���\jw{�!{Z������AX�y�.�0�Jюu	F�|��JF�ji�NB�']����ϵ �����ᥳp�3.�_��C���F Ӏ	����j�WM\w��Ko����z>�N�pO;n��y�b���j�afpP�>Xk��zG.�9*!}z�1���0��x���\��D��F̷&������t���6)tX
Ɖ	?	�R��_��ʏ����V���p�^a�$7���]mq~�������a�&+�EGNB��Ag���V~R����?#��I�+�-8�<'�mM���/|sܷ��IUL��ff��L�^�'K �9[zI�yPol|�tn�Z��׸���~�YS/�����
�s/fp~��q����z�3�W+Gѫ�d#{�q����!F�j��&��a��ǹ�٩>b�!i��n��H��.9�ɪ�YaW������;�rj�޶�K�!5�)�I���/Ut�9G�㋍�� ����>��/�z�՝m^��ZP�hA�d�NO��n�YF�+�(x�Ա+�U�E+I!P�RT���&3�v�Ő�̶CW�`g�;��[�O<k��� R��	���vY�߮o8�Z283�񐣈�oL�����  ��:�R���%G_�d?��g$k�"��Q��nˤ�UIZ�d6�]��`"��u��jW��8���#)�����ެ�xuq�k9W��H��Π��u�=;�t:ǡ�{����S��J���V0�x�V�
P�t>�W�_����;���	��چ���'B,,cx��E��縫�O�pU�:�#�g����B��q�}���|�
�}�k����Z򼋍˪�׫�~�D�o9��7�T���'���+��4h`pqq�h������2L{�$��x��b���G�<W#trz���;	.O3h���<6��)��p���Y�u�&i�4<h�нl�����1�NZ�hh�V����&Rҗ����([Ƴ�b��NNR��0����-A�R{["]�FU�#^^,#P. ��/alx��M��k/N��~j�w���f�0C�( ��e�.EddǾ�'���X�����9�)�o���dP�E)�
o�vx\����;1�U�i��l�MR��h��&KE:��O�����8m;bW�}g�r���C5���:��x1CwKw��T����unzr����/iQm�YR6o�%�g������s����m�|�br��'�)W(�B��z�-@�U��+�WT�O�uZ��#H4_��d��.p�$:哸x����+1�R�R���2�Z�F6��<�@� ���A�=|������:����$erN�;s����a~nǐ���v������O�J�u�0R��}�p̓Rs�S�ȼ��;��U��M����*�-��a�./���.�f9���K��^}����ps|{��|{<������~Ʈ��͋�䄓��Ĳ���xM�X�o����ިa ��߷��Z�:cYo:H����6��Z���mo���\�?�𬿸ݝ��,�z�6zu�.��>09=Y��=���~�=u|���0^������.���~���>L�/®t����R�=ٺBX�y[�ё%ںç�qΩi3�eH�-I��V�?���]��I+�j��+� �/����w�'�ӑ⮙�!�;Ky��Z�k��l�4Z����,��$Z��swX ��Z�d�H����,@x7tI�y1�����q55� &��5���s��np��T&��o.ɴ�KAbr`�ɳ_�: ��q-�r�+b�#�?�}�+�(Q�X61`�rL��6c�n��'Z��+_�e��(�0��
�9��o��#jU�9�o`�I���H:3�g����Kg���-r1�R@M���������)�[�h^��=#B�#"��{����eA�t��|~7	 �Һ|b�H�j��>�C�b��,�]�X�@'�)�	|���s��&+�>���H)%CF������	���A�1�-e�44,	���A`4���zMp�6��F`L=,��L�yc˳�H��.Gf����؎�?�P�s��[톆�f�`��o"��%2�2sJ��0��^�P�v_X��-�ΔW��n��^����r��Ǉ��W���ú��J�G����4��4��	!M�8D�
���Ejll,Q���o��u<�'�#����I�^��;��\1����ܺ���Kt�zo>�����ko>ᆡ�쬜�a��x���ru{��m\A�7݅{^���W�B�F�:Ot�w����Nm���o�<o>���yVw?fds��V�����W�eT�o��x�Gi��ov>k���ʈ���s��s�4�uT[�����-�@[���ע����5�S$P(��H��ww--�w�/|����s�.7����53�˙��A��1���gDS�d�r�~�5Uf�N��֒7�#،X�?��~ ��m;~,�٧���w�����-�hFɼR[�;�Z��2����;��3e�{;a��HE���`w�hi��nWYcJM�������I\
ÊV� ��W]%�����\H����L��$����o۹(3��(]�QL4�u���J;US���D-�'�˔�� �c�(W(R-kQz��:���|���$��M�u.��R�G� O���m;jR<�]�j1ÅIjI3N���4N�c�5�?��5���������k�G$e׺� �Cp�D���.�����Xg�xe�^���̒�m����A���Ԗ��2]��sU���?��Ñ9��	ެ�
�Ly�����(���A6ۏxM��E+�2o'}f͡�5/**�9�
������q9������<%��>;�4�y���ڵ��:��
 �y�o�M�)��U��*�4���a���Ok��Ɲ�I��E�~�x{oT�{�����s!Jj|�o|���H�(}�M�u�>�t��/���S��$U��F�:v�f?�G��%���=I�Lփ�=tm�E|����zRɩ�0�7B� �d~��>ga���8pa(hR�O�QDc�Y�ԅhۋ�G�$˖T.P�$�p #3�ϡ%S�J|t|��9��m��ζ��4̕��a�}w�PP�4}y�26>����i�d�@�lSl�t
JxT�ݩ1t��cԜ�`|�V�Ͷ�CO����ZⓀ����+\�J�4(ԢXx:3m(�N���^�>Ι�9ڑ�n��-ɥ&�Gg�-���Z����>ԁ���о�,P��;���]hS�ǵ2�gOf�	�|����6��'�s�M,RPV����3��/L��z���:������������H
�����sg�bg��t����n��ڜH^~x��ʰ_���y�+pT�h�:���:�m웰��ke6�
��p��m֧MV�A���m��C/�ޠ����|V��!F��P��M�q��ܧ�����[�8���7�V�	�_��_��N2?�'�P(�C��n65ܑ�
;i���V6�ؑ�o���`�k��]���u��w�^����7�#v=X &��t67IIII�]S*n�h�����X�=2W�b̛T�s��Z
��?v{�]�=��P��>
�/v�W����*t.X���Q[$����+��}{��.+���oV	���K"}*m�xص���%0�n1�8Z�ņ"�nn���ϭ1Y!d�F�H=C=���^5��oH'�Aa�C�6��+�?2jG�P~ƪ	�2�����o�m�.�߶��Űi���ױ�<����\�Yw�&���Z+7�ɚN@k�[�E
�Zm&��i�ݿ#�z����x������XV�������4��m�'�������6���(U JL׷x;\�ۻ1��X(���%����J/���a�2�tګ�-�=*�Nl��,�j�̽6�{���Ͽ)e�?��کo괘�����WPVt�y�RR$�) de�g��P���F;^�┢��#N��'������vL�D��W�#�#w���p�dyM9S�un`�sg������B���HY��-/��hY���ޜ|<��]x��rZzV�Y��訄��ޛ1%��gB��Uɷ�R3�^q酾�_eF3�~�7�͛��vj�(������K�b��B���9|�mr���MPF79Ҕ�./i�'Y\a��b���Xa�^Bǁׇ�']��/�r
g\���2�%�2�ο46E��G�V����Le}q��x�d0��#�a�y�����a��"��v[�½���k���l���@m�����}	�`G�F��{�7��5/V�������!��QvDp�V��+l�U"_F3���'��0c�RL	�sd�Fԣ�LVkR�;S秋��<�jj9�B/����N���Vz��y�Q0c�>��w70,������hi��%��[�X�9�1`�9*�u��o%B^��M0�Dp�p2Y�����e���iWp�frZ�yu	dqkh|����*���3��DI�d���6Zr@�oo���Hq�S���bt�FO���E�}��h0Η8�������[n��d��{/V������`�W�\�L�G3�d���
�aln����	t������7��̽��f�i�j	j��6�"��jK�k�Q�˖��WZ�zZL�3��9ҍ���r܀Ɣ�C�`F(�-��x����#~�L�(6/nn�-��C�Dlr�N�ffT?��R���kF�M�� Sf��lOvݘ���Y��g�:��E�-����H�������j�k#Ҁv��iv!nE,	b�[zσ���6� YP�ZI�����;D$<��jV3w䞖�%a���.ahi'�Ћ��fP�i
^��"Ek]��'����So��ut�2y������,����D��dE��N�qfϣ��@�q�� ˌ��e�y�}���u��Rh���K��xH���Ą���֞�9��>#�C�� m⟋8��$^��2�yz�{S���M;���O��j��k|.�jN�����sv7�."�R�-C�-͞��L��U�C0���h�>ɨ^��n6NdW`����ȓ���K��������Ct���aYM�����4���
VG��b��?6Z�e_�������X�i�P����eN�{:�%�5̹��'��zE�.���}:�E���Ff�4���%I��`�՚10��h�>X�������&Kr�Fˁ'��˖iԬ;F�>1�d�26��/|=;�l�M��ڷ5�p/=�?c�(��R��j#�3��7��M4_b�W#���7S�u�_&;_F�D��dkf�h4�D״�{������9����S`���X<�Q�P�訡�r�t
�
�O�E�#QۖG�}V� ��� h�rlb�lq�铲�%�t��zw�o�G��9v2�'tn��]u��Wh=�^����c����kzM�lJj���6�(h�h9�~�u���D++�\5����Ȉ
�*k��%ZW�`٭�5�oT��qA�H�v���]S_����l�r�O���L'�I@�h�ƶv�m�w�tA�R�2�`�"#mC�׵���++���K��N Ѡ�I��ޱ��Yg�,󱉕U���L��E�Q���\ ���r�����LLd�"�9��D.�T-�����K�d�~�ƟX���<�
�u,�]��W!n�*��X�T-�j�(Ǚ�}`;fB��~��[�+�.f��۲V�R��R���EP*��-
΄}�z��0m&C���N�ѡ�8��OS:��|�b�[<��Jn���S6��9:��[����(�+i5��|R>�t���fL���8u�.���p�2�kv#+�>����~$�Q�Vl�j�~����M�YO�.���K-�.Z�X��)mudN�P^�o��v}*��������~g,�P��7jz��|�4�5��&��k�<�4�e6��4������ ��)T�ڄ4Β)L�N�����?��LM�u3�yD�����|�\w\O�ǿ?��<	�5j|#|�_�L�j��O���5�ʓ�3��A�Pn�U�[jj���mOK0I��*��ki#�/F8�[�!-��w_����I5���+Ѯ���Q�`EEG�����$^&�P�쌌B���mmaBK5#�*��Փ��'K��ufc��@���d�ȕ��z)�N��L���}�cwK���Ɲ́���pn!ł�?�'���
��7D9���Xم M(���7K�ta�~�&tz�Ha6��ĕ�:R�3�)#1��[�dfr"�sۨǏ-�> DU|����1ޚ(!O,�j�pw��{�����М�Y�M��>�⑺҉�8�¸P76�q`�Xn�nue��g��<!&���l����H���G�(����j�rs�	!� ��2�cCm9�sL۝	�O��#�����_Q	s��a��Ӈ�U7�XF��ow�ξ�;P�mR
fx��ͱrZ�3�]��_o3Z^z�{���l�~�ϯ�e�V�([|�R�,"QX>J�����Q]�|-P/K�IC�-c
4�������ڑt��D��k��twJ��W�Q�(����ik�+���T�U��; (\t���q�m2�S�hٳ@� A�T*X�P�B���c��I}�X�?�����%?rH�>RA~��.��;��p"��ݣ�9&��-GNth�Q6�C�'����'����F�\da��k o���Ȣd���!�A^\nP`ɸ����+�Jy�(�4�$Q�r�Ӈ�)��ɯ��.o���77﫩xqu�P�ڲT�0��q=
akU�<�th���=St�QN��e�`��?ߺM��
-������0�z*=�8��%���R����V�����i�uq�)i�����+jZŔ�쭣i[�蹀^HSƈ�(����#�������f-O�)�:ml�u�,�jZZZ.�}炨�B����B ��ރ��B��78��_[�.68��O�Z	%��H�5<�p�U�'/��X������#/^�C�Y"L,��
��8%mgE(�U￬�Z�9K	����T��G���.y�=���jPx˲0(xc:c�zBΎ*��_w�`�J� ��~�{`����%ӵ����&���lԃdS"W��G	 �UibZ	AC�_>���+����E�O�=�������>���L��hH�L����O8/�.oe�����i�U��s+�)G����)��̕����Y G�o��)o7��j*�M[/�dʵ��*�4LJ8�M����' �m�4���;�r���Kh���J�u �5��ɨ��e׎�U�e��EE��!����2I�5��1��FklTQ����9n�����x�*V-�����m�,#��?gV���~!>��1?��ϭ�a�_e��mg{'����l�@��>9[)�ۤ��o��j�NUҭ�Rhj䊸��>
�JKr�v�Lh(�ٴn�n�@@xSN���Z_�&aZzzު�yt��My����~]��0�z��r�%��N�;�b(/�m)�zc���'>��iU�$F�G�0(��x�j\ �hMK�>YI&�Fl[AXeo��]�GB�2U���Ļ}�د�4�?�'P���ҵ:�лl��E&,��_h�kx�))+�b����G1�iZ*�c�/|s�.426��s��/�謃q�ϥ����$�$G
����Kׇq�#;��W�<�Ƭ�<~O��#<&} o��ɺ-r�/�1�	�jOO�零T�rmG����+�fg[��'�fKѶ�ՁnK60ˡ����&U39;K��M������Pо��^�!��m��C׀_�j���p��߶T�P���|{�%c�������=���K���lQh�ǭ�UU.O�H�r�91���z�b ��U��$��S�����ExO���C���JNf6zNzW\ϙ�>!���N�W$TPRr� �˔x�on�|ߛ�k!�$L�1]� F*�l/$t�^�{�m�+�;F7�:6U޺�ޞ����g{E�0!|A1O�\X��s,t"����t��>Y�CxW�0�!��1j�II�K��v뵑!��*�i��}�e�~��8��ډ�����c�L֋����T⋰|q+�'���i"t�����>ޓ�P�<ة`e~�'~U���)xZ�{�3�@�5�>�CJ�ֶԅ8]T�����i���,I��Mv�G��0;z.��A׹R�+^�q���	#$<�}�ԘFl��9D�/����S+�Z�^��C��j�ř��&c[տ�hc-�y���-l��&Η���܇��r��Jq���u�6�ܹ���Ւ,=U~���^�Bk�_,Ɓ7�x��C%se?�������y�f�(�l�,u��&u��T:�F��������-��U����':圾� �Ue+�)�0,�n��RVR�z��3�?��}fɡ��ÄS ��q���BO�O���Jؒ�N|�f�;HA��|�Y�%��`k�z�w���������Foyy������R�p@��Cy��X��م�rB{�Q��qз�'D�����8��Ye�����ԛM����b���� �ur���^7v��:��G������❃��V�&�ټ�D}�E��UL�u紉WL���4�U�uv̙n`��N�r��E2.-��ѽ�C�H�)a4W�Q{+��旌����(��a�=D� ��4_���­���>f���������;=	��?�(9�_3�~C��'q�?���$}K��z��WF�Ov|@���:Hߵ��RʙD�hC�4�����f��F{�������]���Y;��>$�'`����d�xWr~�N���	�I�[q��8��ҟ�ܕ�*Jm�|?���VH*Ń��+^���~6^�<��96O.4�<_G(��x�y��ƽ7)���i>��-��E%���Q��z�����J�3W2{�{k��'dp�Ņ�W����h�B�9����\��W���6o���!(�?9«�2�����!�Q����IN� �q4���/�]I�{�eAsg$E�? ��ސxI0HR�0��w|I	ül���|���o���h!z ���-��}5S�9��9F�e:tXC�Ƣ]%�[J	
Lk9�)�>
�G�3鷖q��ae۾~ñ���.��jE7�Ld���#I����3�7^�uLZ:g����%�g�ū;�t�&������bPㄮ H~� �9����X����� (���J,=;�Ֆztϲv��1K$(v��;֫n��n�����뒆J$�nS΋d֝��\*�wd�C���P�ɡ_�xݤ�xݢZ���q՗I��h+�a6h�8h����'.ֶJ����A���is��?ǮH*����瓳�m�zZ]� �j�H�H��`"½��0�g̷n��.�lg������Fa2�������NM�ۧ���
r��&3��c�eqz\cD�Lʖ���8a��MǾ�3'~C�T�� ��!-��'�aq�]}3�B�)^��a�2�x�����a�څ�l�b�a	Խx��Uv��.m/�-�%D$(�.�&���'p&Yung�P߹�<�x��8^־����M�����P��4�Q��H��a�)���E\
��P�	`��H���e��������!h�,էO��r�������c��0�f�4MA^>�x=�dpa�X�[��_eJ�t��W5Q@��h��x��*t��+�i�� �߀�L*�"f��y�h�߈�NdX�^�0�P����
>AARv>v�*ߎ�`�$�C*���L�;ߵJ	�c�)�!���o��?�ӜҰC�"�#ei��X�+��/'�ff���z�ס=�,����p�z�yt�׽Oߜ�bT[~��k$�^�;ڥ�����y8�$0H4�F�g	�$B 4�������ͣc�fxngE�s���t�{��}\�7���f�G�����I��l��^M�sg� ���S�GT�����Ȩj����z$@��� ����7[�#�Z:=+k}Z�l#A����ʑ���;9:(�*��p��9�uܙ;7�-�h7"�����@F��y}�~��k��Ԡ�܏�q�X`���B�,���I*�z��7ݸ�9�������m���4�S'��+����X�� �4Cz�ŀ�[�N�Ή��[�������(^O�+4�x4\�������eo�{ȅ"4�tʰ�KڍM1���P�k��n�Qj�7{�~�N�X�7uJ�o��0����j)�=�,w���t��3��u��z4�Xg�6߼!,$���Q�a��Rz5������9��F�����p���W���4W��99µ~�G[C	��$8��[o �E�-5!AsΣ'�bCb>���.��%К��Fn�o�1�Q�é�����.���I�&�֔W>��9��mW��e�-��Z���O�M�k>I��ϰ@By��v'\W��Z)�<�"-r���Z��'N�ИՅb͉�X�<8v�l���2�q��g #��Ԫ�y>!޵���#�_卲5�D ��=��XE㟑V� :��%���S�[��7���p��8����5K�i�l֦�)��h���l&�dxKCKK��Z�^���v|\�A(�8�����>�*���x��l�+kS^�D�6F*t�4/�+!�a���-�OfD"�����෻�&>>��9��k'���Y��K�<�B������I�[��{�2���H�=\ndת�R�[,�*S-���g�'y5���Nj���P�v	.�o��1�l�c����0�ֆ�j��q�����o�\�'��`z&�t�i@.^9�)Nh���4�d䣽%1�P�����;S*�VBE_����`�H?>/�-O米��*!Ў���~�NE�,�a>?���Ͼ}.Eߣ?2�0�?f^SБ`���-}�oH
����:�
P-G76�c�kQ}�$IUy�X��C�V?{~ȫ`.�'�xhl4>���c�������2)m�/{M����W�u���2�o7<  ��V��o_S��3��;��1�%����-��_(Y��٪)-M�_�G��"{gϽs�Sz�|B�9�P���g��cT��@�г��.�![��S̓-���g9��񱚆�ގ����V�Ý�����4��ic��[�t� 36�r�;y�#���O{��i�Zڰ� �3ҔS�(M���Gʑ�

������/��L�m!vО��Wo�W3k�*�qq���|���#+����gw.Z�R`R"ƺ����z������螟���#q2���٩�ަ�n\-�+j�RZ:9���$TTV���%�/mj��R�:��3�F(ޠ��~J/6?��Y~�O���	�8ȸ
�
�F��Z�oŭ^�P�ft��ʛaB��Eq
^�����2D���2���1DO{�0:��Ꭰ׽w4�J�E�Q��}Q�1~>�����Д���m��j�x�S����7s!S��	��k�Yϊޥ���/Ü7Ajύ����?��_W�ɩ��v���J�G�xj
~�(������a��������S\k�<�Ш��`O�׈��7��MT�<�%w��p/��؛O�̥�!�ul;y����.?�gIgPK�8uN�1&��L�)��Q�r���	i@�#�,-�傢b��)��u��K��9��όz�\����GnB�t^�ӔTSs�j����O/f+���?iq��_�hvX3b�������w	�í�4��>�?�����k�->�@e����3�����v���=mcd�a��`�ڷ�q�P���3��9�Z���.��W��p}Z�+�q�����M��{;՘V����h�t�r]���(=��yo��8��3�b�Mpj�:�p5���7|��F��T���eī�d��AF	�����=�6)4��F�ع��^������ăЖ.���p&I�l�����l�������[l�3k@�`�? ٿ����7��{ǒ��O
�#َO��go:&WT�c��{#�wR��B��)Ć77}B�����P�9��
Q7dT�+���{w
1�Y��C�WŶd9�ğ�<�-.�p��M�M�'�@i&���62�߈(�[�C�$��c�>� ~���!�����T��"c7�'��YA���0���M5TX6�H�~�a�( wƓ���%��3�4y%���C}$���l�uƊ��?1����4k��h̵�-d��}�|K��.�Z<�d����R�P��㵶\���o\T�>�����Y�_�&�������w)\^�#�(�t��C	�[�e��6|X��ى09]��-ԲQ���c�u_d���	�Ա���_�2��Hp��r��l,.ˢ�ӈ�.����Ood���ƪ�&���(����m���>��\M٤�F��b�����cyd����^���-�'/��a��vA'����ٶ�'4���I97C}=��Y�Χ)g�'���ြ�O����	�p���w�ea$�NW^�"���5��|�fZ���md��B�ү6xfV�`�-*�C�歒��8`Ɲ�'���c��vH!�E�NkU��TH���fn73�&�
�&�^���ʔh�0r�
�|6�_�5]�8���]����>�~n�D�
�Ҳ���>�9���7�Z��tx�5�O�m�76�/~W��7=>�H�\.�C�9�uּp8.O�N��o��������vw�I��d"����u9��s�����I��c��@J8������o� Y1�2-����*(��fHZx�����$�CgU��B���Ch�L�ҫR���5�O2l1Up�3/�XzC�O�����om�������/�J�7|�<�<%uIs��o�U�yC45h����:�닖�?7s�v����~�s$�j|'Y+��/�%F�H7��۝�2�d|�lM<�<�0P�.s��y�-ŉP�͑A� ��dT� au��!U��oj������J�f� ln�a� ��j�o�%����4���2��\t�3Y�z���]D�7c�2J�y��(��g[�ͤ���[-ځL�t��1I�����0o��/j#:�Ɠ�a���q�i�12|��,���?~�R��S��As��Е����k�O���K�����{���I�,nC���X;N(cɬ'V��f<�j�����e�������"K6�P���?e�+��=�9O��� �l�ܭ��?�cc�P����ɛ>>\�:1�����z���n`��w¹�r���{�]+v��������*[`$:�$�p�s���͠���� ��y�#�cU4w���+8��ٌ��Ӳ�7�9��]V=`��')1
m� �:N����i��ێ9�������J�֛�ߜ|\)�14,X;�	�h�Ը��9�>;��`iYY��n˭��R0ө?����ZWW�؀E�%�KuPP^~�|ʉ������eb�4J��~H�%�tJ|22~4rL2Ӥ���V=�2��ƴ��ӏu�������`�aT:-���|^]���b~�A�lT�H�k �~k�Ŧ�>~�!V4>|D��Ǜ��@0�P�S�5�h���.g�j�<
�IY<p۸y�����(�	��-B���9���M���ݩM-(�2�����#�OyCelhii	�2����j�	���%5-=��W�װ�_���5��*��� o�52��%GS3�N��Ǜ0>{�������>��c�l8��a��w���zl]��X����!"2+�|<���h�7��`lG�r��_w���23xܲ�1`��P��1tb���gaߵ���sa�ݴjbb�:�h�Z����с�Ց��R�����c*0`M��P�x���{ʤ'�����-�m��e�51�M>���XK-�b]�e	x���kKK[������F�D�e����jee�>��t�����1�x�Z���w�~��#�}�Mm�>�:�
R#���I���bA������m�%-m9�@�Pk��=��TK���+�ԣ(��)��{Qz�ZHC��©*/g�.Ѡ�5^�kq{��������O͠�����A��ZZZ���Y�_sv}@��\'��?(!)w?�g�Է�O��$}���2��/��Aa~�����T̝fty�� �SM�K�����^D��%�?�bq����g�ٮD�4�T����������y�H:�+����(�Ȟ!c���x��+Tq=:/��uk�
�%_�5�Î��{M'l�L����ǽ�|�`gr��Y��`!ߞ_�����8�����c��t���Z�G++.��GOa��W4� L�3��-���?#F�+zM�(މ-t�ږ�>�
��"�Vm|�)a�Gň?�-S���<L=���?9c�Ţ�z?����L���U����A@�鸖��"��"	O��z�iJ\:W6�h�u9��U�K�K;�`.��7G��WT��SV�V·L���������0ၞGn�Tُ
	��Sv��'�1����	��;�}SpG���>�m�L�����jIѢ�vɠ�I�ņ��·��
�F��I*�:M≴�� +�r�*�p���7���1y��S
��a�%�}���o�'�T��F��;����z�2������	�)�7�MP�?�V�1k������o�]!S�d��Nۓ��=eWZ��R��,<���!�T�G��*󎽃L�*7�f��[/�v�:,�'� W��'v��Z�1@q���4K�"&/槰p�O���l���==N0��B^z�M9���W2���5'���%a��q���2�U�z�̤�����k\����̙���Q��K����_�d��*7N;��O]��YۺV�h?����>".}//f���1�4�'�5�/�'w%	Ӿ.!I�ƪ�`������z7��k2l��|LT��d@c/xi��#SA�(�Ǧ]Z�y'Ȃ��׽PxNQ��4���������V�w	v����d	���T�O��W �i����1��O�|b?�5�z	K�{:�&�7n�)z��}*�5c35�t�X���x7�Tt�J]Eb��vAKy6�$O������R%��î\��,拑
6�3/8���H�?pJ���>�I�U��/c;�ߝ��v��r0�R��B�qo��JuQ��]M��V����{L�O�����?N��N�0%lOF�N.�5�o�1w���x\���Y������-�dK6��n'��w�<@N59��;N5�{�o	#�+Z�s�|b�j�k�4�����$·��!�,�9<h�-\�1��x�
��@�R<��\^���a�I\�l�)��g�̣���n�������YT�Ǘ��z�+��+�ƭ�C&�*Se�M��j�ө;i�앲A����?�R���꘳a����(��U��#�������T�n�`} ���L�Z�8����
"����W�$-�R����/T��|����?�nf�?w��}Y����q�ޘ�x�ER���f/��B�^�l)2T�`���Yt��h�X�Z�q1�,-D]��m�иF(I��Q����#Z�k6;�T3赪�}�1�����2��U/� �f�YH=;��݈w۝�_?�QL-+V6'&ǄM��?��W�ּ����?XۇR��8r�Wvef�R?t�iw�i>����!:j�6��+|�������/�����uܓ&RK�*��O͇{���x���e��WT������7u����}�_���+�U����s,f��ƅ�ݟXo��{i��b*�����gv��f�8�AȷV�rA5��~�;%������ ��!~h�-,��;�T����U���#L��c�Z�t_ Z������.0�,P���$V�J/�dbtlp��i&���Xa��(c��{�ǽ.���6`m�R�t=�^���e5�)2��g)�K z[�����2��9^t�KO���I��c��i�|�a�q6d�OLW��ah�j�i����2�� ��t7&f�!:m㒵�(7"����	�/0� İ��v�� -���w3 G%sL���a��ۃ�R4)��V��fs0iX-����f�	F�̚V�-5c�5{���;�+I��@�8&�j�ky������/)�/���oD�&��;�7wG2��Y���P�k�F��񕁉
�7
�}y��!0�L3j/^�a�1��3�:G4mcI/���%�xQ�=
�Z ݳ�2��Q�H�\�U��*��r�#��Ɓ���	�{n��.|��M@�m7�l��͡$.��		��Y��E��6*�ZO䘭u((*��H�M�[�l��b�-4��-�������M;��m��a:��(�*H�M����10���/���A_Q��d��݉�?6�[zș9���N�
(7�,--czYIv�U�;"'� ǘ�9n�^�����F�tk����ņ Q��)�A�^���5��3�5��w��'������p��}��a哑S��U�`-�S��̭�{"e=�@}R�Z��f3��UT����]�q�Q'���V/V{�}S�(f�C��Z)���I�?j� ;��\2 ��hl��P��W�`��3f*�+���ppZOX-��%�ÿ�9eօK$|���i�h�7e	|�yЧ�f�YuQ n�g|�3�^CI����Cs�O ��j��5�sOjܕ. �j0��֏�N��N�<����,]��r�kV;�p �U�j�NS��8�ȶ��?{�j֬}��0���T��0\���K���4_��fo��\m�]��L61>y�w�2
�;�v��aN��'R,A��w����G�L`�k`H��ï�x����QI��DQ9����t�6Uɶ����=��w݅v��	H�F��)V>�8��
P��eC���c�Rm>NA�Qu<i{�� ѳ��xYFǳn���ߛ����"�{��RS�؏�2�0IMʂ_�r����%�)2��5���ǳq&�	�	&i����N��L s�L��L����Qi<\���R{�>F
E�����[|����Al�Z�I��������(���J���@r��oY���e�M?��Ş*��c��f�.ں����\�yӄ���vR�:���=H��a;�+)n��_��Wtޝ��_&��#����=�!�#�2!�n�)\����΍x�3���)$����V�d��VW�ˇM�Ge�[굖{�絉�3�K�l��9cI��A�A}##�h�e�[p/��l������B�Y����)Rr��� ��ԔL��ղ���غ�	��$�����������'P����k��M�~sj�� 6�����[Nk��H:$�|��lʧϟ�����>��9611�׽�_�5~�s�k�{}���a7�$DcglX]�����ctu�%���囟R����k;(c%{J��'��qyGț)�Ӗ�Z��Wz��Yx�2����r�ir_^0�$�%�X&��@��L_��/ʌ������~�)��Ry]Aycd�O�4�ݿ
���I��-�b��!D`�u}���KV��׿���`���O����/C�5o�A�P�S����'{���f	��m^C%��i�j��S�L��g	q����<(���
#������Uc��vYe�~����[����8��	Ӷ�Ь�-��8��v�ǯvjЃ"�/F�Vd�@Q':v�X��l��l�뱚>">Z�������"}��J}z����f#ڷI�T��J��c�B�w�wqC����%�q`е�B��f�6�'�x^�~�G��Vkc�W�u�f���磜�DO$���{�"=m&�z]������ �HTq�Kl��2�x�V�S�(��,�Zj':8Q+��sK���d��>A�)O��RS����B�"�a#ޖ�����Xy�~S�������ߕ����Y f� ��\���F=��]��jJY|#Tq�}	T�G�����5� 0r^^YQ���~�:X�\�>��"߳F��Z^����9nu���MC���:�(�����v-�����g���Q�E9j;WZ:|��~�1*�����Q�������gN3KЧ��x���&�)��I��RUP������eB�*����,a���ˏ�����]-�����
f��U#�+B-픛�b��A������Y;����T�~�����pqީ�˛�U��#��)ڸ�I��ɽ�W]�_hoD����eeL��}�ā�b���+�P�ti��4ѪR�{^@[h�,ţh*��K�&���޻����eJE\�P�I����I�$��,n�m熍*�c�n����M<A|�X`�K��]�����ƈ���4��n�$ �mēE"6Z�xR2�����L!J��.Lg�E�x�v�M7��R�'H)	F���ȯv��J*��xZ��s7|���|��g��x���X�6cJ=�����:[�����܉�jh*�<��?�f��[��5
��>�0DΆQ�L����w���R}��`.���n�v�Bk�x�K�ڹ`>=#�����8O,X[,*��P2�?���^���&���:�~ ��!'�z�KM��n�&��t�(�lF,Ό(��tp�����R�9�-�����N��)��ε��y��C�;���Ȍ=���UɅ�/�s��-uߝ?=3��B����
D����ũ�_��wF�Z��G7����՟�*����zƿS���>6�'P3U���h��.}��J�Lg��?�G����L�5�G���K\)��Oҳ*��ʤĆ�񠻟��*K��u��q�g�$�b�l�#_22�f*<�&�.�5U 01�$zЮmj0+��̇�H��~�$�^�C�"�6��ī��Ͽ0����� �E�x�Z	U��+���=)���ֳ5_�����B�B^��Yht����I|�%p����y�XYE9U�7�8y���×��Qi;2�_b�	���	��?��:�����_B�P$�C�k�" !�FF�%��K��H�to��c4�]����?�zݻ{�s��s�y>�������<G!4�@�a��A�iO��D����������2���D×}Ԗ���}3�PS���k����m�y˽]�}�O����}�K�I>�2���SU��@al�s�S��Њ�����F��Dw��z#!�m�7'��\����&�WU[ϑ%��-�T��㠦����I�f�,����C��d���]���N"�KgvS����X���H}�^��K�=�ěq?HwZؚmw�:�� <��$�ᐽ�UU�̫����j�ITS9fd��)(k1�@p�U�*������E"P [��5z"��[��_����e�}ϸQ����II3H5I'$p>�<��9���K؂�2��p��I&Oqy��1����Sz���o�b�������vs$��!&"NOFk�a!�m3�S�UZB�5�޻f#�#�Q�O���H�_:����M��,X{e�'�uMF闼��e��*9�X���r|'������$T��q.��H�^֧�5��[����pw �}����?5^��'��/�4^[U�'�k�uϹ�G'�͐E��Feվ�=�Bl�ӟ-̟d޲d�S�dn��7~�� ������-��L�	KN���vTm,�ZT��6}`��@l����\�M�ndK����蹹C��MKTo���h�g^A���N��֪�mO�2�_]����M:a��l��������pg���Q,_V`���� �S��^�v^��w����������d����a��y�n�9$q9e/��6��J��Š�; 'Kh�����T���vr%>����S�S�/,�?'hs�|��\�E
��&#�$��l���-O��y��4�G	��ʕ��[MN�3��B�V`P�NY��Y���:�4��!��B��3)Щz�'*
E�V�X�A�߫T<�5�7�P�bŖ�	���_ez&���ˮ�������\S3{��χ�＋��]G�ΟI5:-(V�lޛ*]m�����9�]?<SI���K��<��N�馾��G��lX���#�d�9��?�(����6�_�'�WH�;�vR�w�jJ�T��:��]]�qR�{p�XMIT)7���0*޶ͳ��y�l1�˪8K��%��:"}���A��U]Iaw�������[�=�˟���&(�}��`?w�I�L�O��N�ф7|��Ӹm��Ϥ$�P����x>�+M=�ϻ��J3��땫m7�h�q��W�x��#1=]��#ƾ�Ga�E۳���/ň�{=lm�U37�Ǖ�f�ܩ�������*_%�p�n�>?X@���llk��_^.s�m��X� #b��H~q��|'����������r�f��f�����EEp;����]���\�}���ꔪ��Bq��C*�7S��3��]]�ە	٩����U�����pR��)�+�!�$��N����X�(����0GT��Q�*_�0�7`�� A{�Q����yZ?(���3������̈�G���eB	�e�@�PyB�ބ��wK��l��B�9z�KG�^�[om��(OfV��r�c&W����jps)����4���̅�#��w\���i�C��\Y0��#c�~z��aa�X}��V�P}d���8�Xϯ���o��?/���]�D�(����T�Ȩ���`2Q�V�Ro*:0�"x�<i[~�G�q|����/�dtcgrrR�Q)9��}|�\Ӡ���k��^��D.�9�fYܸc=A/��v���&�kd$G���tf״po��	�C߭���g��(���͵gT@�Q-��G_I�8%�'�����A�m�{��n��6s�I����%s�/��u]7��Q�����ѽ5S�U������r���_{�i]���ۗR�ZD
�ŗf������-f��?���=�\u��3j�|l0?��CU��������Ө��w`i����X
�ppQ�Y���se�s�S�BV^~-$
�&''q�lKQɔ����-F��������?b��JeSf�n�������<��h���x:P�`���z�y_F!�@�Z�)4լͣ�(�J�4���	_){W���r����
�Gt��j�}J.����{�Y�\ɓ���������'AfY������r�|B1�?���@/uȶoQ�)OOa���D`�`䠖����Ces1���AȮI��;���IL�Ū��ģ���Cvl3V��GFF�� ��Z8�	j|���ztĝ�{Y�u�"߄��T��
�$�E�1��3ssnh�T\R��w#��C���hd����c�!"<��.6"���穪2*v��|����M<�z�P�o��S�[y"��i93e3����wS��S��,��jq�OhgT��~���Ԗ�N�|1�
�1�y��y��a9}��������>�[m����Ԩ�pO�͛�"g)����Y�=�aÊ��*�:_�"����aۃ�i��R�#z��d���PZX�5C��s�J<=���CϖW�������ܛ&:b;�y�B�:�pDZ�Q,'����������͆i���,�G�0��Є�f�{�<ƫ4Ct���|�.ҭ����WBh�����Qň�/��41���Q�����/��=E]�.	8S9�IkԋYm&�:���&����7�yN|>��60�h��%��.�X(��~ҝ��Z�LvN~q�X��������E��7#�rڜZe�N <�O�_����9��}�}�b�_*����#܂u�ށ�M3�+�!F^K���=	����}¢H���XlП͘���4����$��T��k��m|a���oEzH�!���oV�A�;!x�ԩ��B�*�m��n�V}��=����3���EY��-isa�y�;O��[�Be�5���d�
ee�1�D�n���m���>��Ƶ��@��k:�P��G=�J&+�2�
Ida���<i)�'��,N���Tl�v}ҕ���;'u�
��"��� .G�$@�˃[�������m{[7%g��;���:ipz���),���f{�bj"���Z��	��,�n��A�˱c:{L�\�����|��: f��p�f���#���6���i�댑*�lH%���W*��V��J�c�3&�}~4T�KU Ff����)ʒ���>��ږŷ����	
0L"�܆��D�*�j��"�+�`��$��27'^��C�V��0��p�u^��L�Ք�b����y}f���hrR�q�17�6?��=Ȟ>\^Y�'"N�j�i�OHX^��DZ?���	�laqӯq��t�~7�+�](3Y7���d��-�E��*���?4��+��54����)f��n���m�KU�)�s䓑�ά�a��;Hk'5S��0���b]w?������e11����>4�i����
�8�'�&��V��LZ;:ƈ�G}��LO��N�c���-]J3�u�m��N�A��A��4�;� �E���-7M�[�2/���5�>'�	5+�fs�)���7�"�G��Ta�OV�㹾jN�ǮɊ�GMB��&�AeL���{��(O����sq'���=Ҕ�H�8���敖v叟}�w;U���^�����v].�%�'��C�oKfl6Gĳ��TG4&_��[-�~��$���.f�5_H�~ߢ�>�Rs����m0''O��E~�6���/��`I�f�
�RPP��Ԏ��(M�ڛoHScOw8m��R����d��i��B�G�g*,��HF��Hqqq���>rA�7�x�a(��*2���m��a<���ͷ��w��6�]^\�o��fc��ST�|��F�W�-,r�M`}�̚z��i55�R3m�IPS镌���|Ysj`�LfF�����dH`g�x8ߓ̜�z��T݉}0G�����LA��?�:w��D�9�)���\���=C�!C.I�:�N�N���>�q?E�����,��:������̛>hsR�S4�Q1��k*�\y=g�}�d�o�D;�dL�8z������@��"���� \�K��4>���mLK���b�p�Ikx�U:�_}Љ�F�xq��s&ΧΞ��F|��r���shs���d*��%:1�9R~Q�����4D׶v�{�-k����wN��M@ގ��Um�O:P����Sȏ�)G���xp�ۂ�����\mcn��Q�y��M�eqIa��;�A��Nx������i0���v���+'KS��j�����)^ؿw����	B�n���aT�����H��@��JR�YZ�[�!��g�E���ע]�<ݠ4��}fL�������ޙ?�[>f\�s�����k��Y�kU��8�mI�ՙW'z��rH��*��Sށem5AL�������>mi_�S�_���w/P��U�\H��3XJi"�k���� ��C!Im���Fg5��XBj
&�@V=W�pދ����8������}R~Y�.��%w�2��̪��np)�U��ժ[aЩ���to�M_8�$���w��ӎ��ܐ���t̫�Yפ e#p��U�����#C�$�]��\�����a�1mQz9I&S��6�xڬ���O<t�u��������B_�� Q���С��ޱ���R����2���\4�rg%!~�G�Gn-].b�36x��=z<CT/&�M5�c3?rF�z@��G�`�Q88#;��)�)ܳ4eX,3X�:[\�t��m5��ۖ�G�%R
��������ǊN =~j�����O�l>��7��'rQ�ym��_�����9� ]�x3�yyVNV�P_BK0L����2�ްA�����Dϐ�	����#�����ֺ�:��3%�����"UUՉ=����|��;�Y�n]�Z)@ni�T�d��3�I��/����TWG��_����<���J�)�Q��&")8�&�$!!���Sn�)����jd7o��F�*�O�_	n�za�&G��8�zU�d	�|Q"[���S][�I���z���z�U����ѯ�.�^��!1����+z5p�k<w`D�.����brbx�R�ϥN��^%c�%ϱ��#�Jw����_��f�/��l�Aqb����M���mj�עKn�Wc�W	ht'&�����b:�����4�9���|f$���JxC<}_GaK�ݘB��1=��s,�D���_%���8�o� N刍j�5��Ҩ��2lb�,(�!_[���/t��! ]� �<S�UѺ���O�L �Wѡ��]�`NK �U�;U<�(@V^^��rR嶏��Y�S�):�'d߷�;��6/���?�+F|�C}�"����z�q��{����X�#��%;�RmR��#��Ö̥�)9Z���)}9%9�з�J� 3�Y��A�·D�8K �{�h�)���z�Ø6 �B?V[���~�h�?�ꨰ�Tv�+�͚���FM�����Y5�쇣i��ȗ<� �N�⨱�V����{��e�_�/�� ~�������`k� �T|�`ƴ�I��;�~>� � �.���9U��Ȕ��� q}�Ȓ�w��xoS�9��]I!0��P!Z�<| W�P�f����6��T��5,��Kfh��W4�Fی��O�`�{&�+��=���#�����K78ɛE�*S&�r�d�9��%����?Tv|��s�"�j�e�P?�T��o�U�m+�B>�E�L�z�I=�pV�:<S3T-��<:�G�6�I�?�2zL�f�ۂ� �%"-��̡I.g�
+�rWŮ1)~9y�n��(�?��f����[���3o��~q&r��%)�ٽ�hR���cb��?*'���G����f�����I��&p2ʯ���mÓ��j��E��G����$ʲ��S_c.��D������W�|>a��}؍'�{����񱺇�";ǧB�����7�M�.�Ɋ�`����K�#	��*��E()�����(��3���Ag����(� ���k�Q�:em�k'�c���[�w~	'�W�$��.��ػXT�p�R�C}�:�7�=t�m'�'N�����i�"��� �Ew?��	=B*����;T5�s��V�M���%??-q�Ϩ����R g��SӒ�6�nuUN�ign�[��Z�&W��-}}WǙ�w�0����ё��R����l�#S�I�G��̘1���_w�����l�w�`i�͍��Q���C�N�G�>O-��z�7�[��~�,.�b�o���.��%&>�� @2�Sl�r�y;���7�BBWY�@K��`r�/��Bw�C���985�E6?	���5"�`�]�����#���M�+�$f<��j����"�����<p�[X ��<��٭������� g��Ѽ��k��#�J���Ӗ�+�"�x��э�8��붅�޶��D�~�[��	�ʆ��CV����Ֆx�&T�C�i��J�I����
��޸�K�/�͎��.��eo��W�z�0���#Ĕ]����tdCks�R��_��_9-xA��q��B"���+&���͑{����Id����|)�K��X����$ ǣ
��k��+��hV�<��hhSK�e݇l��g)"�5����&��i!�>��Цӓ�o.��i�K��xg�m��yt�����w�<��i���T��R�"ѕ(��<BjI05ӵ��w�}�y���٪�}�-�|�j&M $�Ȣx����+K���y%����ٶ�]�G��O�UO��d�u�WTsL|�jq�eC�_;�Fn�I�j3�
��E��Z�������=�}Ա�Q�f_���85�)��AE��p:��r���I̟�̬��g6[2���	�vi��=Aҙ�/�3v�����ms�`
1*�E��^f�iz�o!d�*��H��_{�,\M���;�/�K��FM��5v�Y���.����K�k-�������M��N�ll��j�uACΊ����Fm7��o�d
be\�}[��j���1Φ[���	�z��{2���v�E���dt���y;b+����˗�{WuR痖BYO��Vgk
����a�=�?k�P�y��Q�:����j\�Ī<�#��̽��Tk���,���W������ޏ�d���O�қ�4�Ud$תju��yB�JZ��A��l��?O7L$Ҭ�������Сd������\i�vF��@% 5q#��(�Z���(�l�f�֊����m�&Y�t�_�B}=�ֽ�#�K�CH!n�`�_��񺏝oB�����>e����T`�Ϳ��L���C��?�?d_}��)�m���Ħ�
h��p����v����J�w�gp3����b�
���g�GC�QwK ¿W�0�|��;��SE���<�m)�b���$�a5�	5G�'��:�����oT�����l�z�z��.!�ʳ����Ph��\W	��}K0���w]�N�D5����\Blb��F}z�7���}��3���#�&[.�k�J���$xoe;hu-�����-���}������Uu�U	�X��'"�}�$���Y�EfM��0kԺ���m@S�N�.Gzȋ��|�Џ�鼣t�"M{]?��k\����^��+@M����9}����ظ�|	�@ݽ��5���)����۟�z׀詓G�\���/n��5�'K��6�X'�
���ȫ8��IK�zΘ�OD��R?�ܛ������9���'��f��_ݚ{��^/�DC��{m�w>�2�Bc��� l����q��+�g6
5D����t�ht�5A(�$x!f�U��%A�/�XB�dC��8eM��I.�J\���1?��4����v�tw\h�u�340�Ud֩��c�Un]����S����*�џ��2�k9��F����G�K-�yK��O�_����noe���E;b��G���yR��ǖNE�<3;�y�`@ɈCNN���͸��C[=��.�w���6�̯�����}��l����7�X~X�!��ش�B�4��FRq��9A1�=|9ҏeS������x����_����8�G֨�5�L�@�z�GN��Å���������yxi3uM| ��>a���x��<����n��Y��ie$t8D�ea�>}�=H����7�
K;�Dfe�x�
�RmN��� 0j�h'IZ��r;X�[��r����R����wGЭ�*�*�u�� 
'�|���Qѥ��#ٳu
�f��uBڛb����P��l@2�Ǎƥ��'��|�쁾y�s�ثp��,8Y�4�olZB��`��nu�4�<�R��1�(z.�nx�e��2��PO�
o�/�a��j�^���Q���	f�����ۥ����\��*���ovZ�(,�Ƞk�1{�杬����V�<���ˆKd>f��Y#余���u�5�ԫ&�����?e����1:���{��y=#�T�v�W�Y!��?Q�uU��z	S��!C������.<hW��C����(�W-�����0�Z��<�� �r����ʣ�� ���8�˿������n�+��~8Ӣ�>jE�c0ummm�K�'.X!xuEs��d�u:���1�T'���6S��X�Aib�@������`ܽ�{#��Vx�����8\�S�H����K5��O.8_xu��j��
5s���M�u������'���4�MD�`�-��B��z�3/�`��W�>�/禀��e�ɴ��f=���1��A��Հ�a��q�P�(m@�͠�9�����}{�g���?�Ce��aq�Tp������	>9��\����G^m�[#�C��,'�&�7�"���vO����Y�x�E��>�����0 �T���>X�vf� ~�����pQ��%(.޿��7��\���# @��@���۩Uׁ+�Ǽ�kn�ST_���$�I��@���ҷD=��J�Zrdj�U�y2P�ݡ�c��R�9���F@3���c���`*^U1���� ���#��4i.#��?�H��3Kk/GX��0�4\���J]�i�<ƙ�����i�HFgi��vs垢�h����)�C�>;@��K����WVV�]�$1oU�v�V�X���҉;��.G��%���6?u�TU��7��O�M�/�,�jĽ"̑�	��ad�&��؜T�d_����^�l��p�F��h���^|����
��������f�Cy%��Z4�*�G���.s�u�7k4��>o_%���{Ff��4̍i`~���R�m Ƨ����O�f��V��n��
 S�)�06�Â=08�-�;��M]�~*�j;�,���W,��UUU� ϼo�`�z�����f��J����}|�E?�᯽0���o�+I(S���] ������ٔ���7u��x�Ɍ���N�z��X.L���U�j�8~-�3?���yCr�`��6�a�����2�r����폌�%��|z��IkF���'��zGw7v���(�q���]��8�-~�}f^�2�1��Y5�}ٍ�sS��o���I�7�{��-4��s�v��$� ��E��OZz��tT����sB�\�*2������Qz���@'�}��aR#_�͓{��'gP�JW1��`�0�a�=��f����W#��}yrAx8)\�D��t3��\q���3�j�m������7]^�h��&�c�X�����y��j)d��}��}|G�6v�
v!٣:~c�;��|�B��/h�S�|���d/�!�D�a�;����u��.wla��\��"nL+;��`1���Ԉj�����������^��X� �����P�����!J]�# Ӹr�Es�F��v����c�����<v�~J��n���N���}���H��;���"].�J�T�_�pkk��V.de�Ζ�`�[M
Ƥ��\��?��iܷ�JҫFb����ѝq���~p��<��U~Js�B]tH0!�N�e�҃.�}�O������/��Ӝ�h:�d�hĴ����Z�FFF*r��c��du�F�:�����w��2�
�U:�����Ͽ.ͯ�It}}I2���@<�J����؅�X�N��E���`A70Ϫ������+�`	��:o\�q��\��RSɩj�m���Zj~��A��3��ܡSG�mc`v���z�a�
cXusB@'�D���a�Ժ/b�Sr1s�����d.y`�X1"J��cb곜�>?����]�$r!�$��rо��a6��Lk;[��D���qd�� W&�s02��{q�n��Ӥ*b��y��I���W�Y͏x=Z~�58Ew�3:-k>g����KK�V;b��+:q����3����N�$��}�
�:!�/��-@������1��!�Z���$�H����:gL��H�e���8o@	��������a��F;�D1�U��P�8%��X.�wd�ޢL�v$y�i]n�C�ZB�l���m���Jw�}����K,_�n��l���DI���H	�	
�x�����O���x����N��z�G j�c�i�����X��%\M/}���l׳B�-��5N�zA3Z=��y��*
ep���k��_P{�I'=]� ��K�k77Q����~B��%���K��1i�`2[�v�_fNF׉1��p��"�C�����?�������E4:yƹ�S����;��G!J�J�	R�2;�XZoZs5-��Ԑ�����l�1َ-�r�R���K�*��GȒo��ƝW�82��9�b��{���s׷2떖7
��ؤ�G۝��m�]��0�~��zA��*>3�$r�4��E���b$:�|�VT2���Ʀ`ClBj�D�L�ػc�Ļ�~��C�#^�N��z`���[�NMy���r%k���쓵�j=��ye~�R������8Ev����O�(�d!&UArO`��1bq��������;87c��� ���rK��?aI��:4�[��mѝ���~�>6���g+�ͫ��*L���W�"�:1~�^71_W�9u����q
=|?&�s�~��S��� �hIq1�I�m���
�ÔF�M�4�u���0hӍ�4Wۀ.�FH�잙�����i����m��S���sq�:�ɭ�����ʙo�Bh`懄��_':7o�ڟ��(��K�D���,w�9>|-�YN�""w@r|��Y�.��hTB��eo�l��#���)$.L K����`�ug��1�'��3�:��ܥ�Qȅ�R��lϬZv+7�$QF̅�G��� �#���m�Ur ~����d��&�sf7��/{U�&���+sno��=F��
/A����BTb^�� ��C�I�HCC5.}��"����8�*v
A������;/�0kˈ{#�$+�� gY
|�b��-:��j�)�x��f�x�.���t��,�d�����#m�r<�������������S�)z	>�I{^�� ��>)॓t���jX��=y�8����fde]8�]� #�3R�e��\�5����"�����ԡ�-�Rqn�:{�ʳ�1E�7{y��D���{A��r�4K;N�q[?&&LP��|�zK�ݥR�E�w~�i?MP7K���<H������8x������~�yE�o�>�Qt<��e���ҍ8��Qg���:���(�򡰩ho-�j%��jy�
�ޓ�������+�e�[�'�6���$���dE��U
�B�<�F� �����{#��x�_�Q��3����9��N2{TFF�F�!�Ġ����$��� 4��x*���#�I�Ʊ�x��K���[�$�|Q�X�}�Ʉ�����A����g>��3�2
t~�Ϊ���Q[SV.���g�*g�q����k,��ig����S7������KW�@:�c�U2?����>m�:�m�{F+�m+��:�l�/|�����@{�e�s��=�J�Z������C_p1�.�I�"G86_%����?��
��5��5�(��t��	ɭ`����� ���\��tJd�h�ˇ*�#K^��';���܁����A`7���~D���vv�n�)}������ÉB��!��O�:/T��4�d�v)�^��X�I�QI}�2Â�*�r��>��j?��B��} l��r{ј�F�M���J���Eb��xN�wҸG�Fi��v�/��者�i���8Uxu�0~0���N*����7�׋J�������qg�e�I¼��&�*((x�t�;q���ta�jz6]e���R"�k�qW������,Ƀ�w�5��c/������F'K$'�G�6�7�b�L1A�Eq�&�i��+��é��We��j�v�o+�(��dzqq1�B��11�g\�� v�6-�8�l�Zr�%+���H--z@s-��P}�r?�Pٟ\3�	�0��ʭL�ff��B#}������Z������WWWv�a��5g)C��s����st�� i\����	*��YƻcStٲ3�c�f��lIβy3�Ԛ�J�9Ls>Z����4b�+��Rg���f�m�x^�X��f���XG0�<{�B.��~Uk>Z��8l'݌�$�&�#|��Puw۰���c/��H�by��<�{؍��U;%L���� �Z;����������R�q�"���}�2]�r1�t}}<}P?�L���[�N�s�$f����jc����++t�i�igș���󉋲�}{,��I&���Z�]%��O�q��Ѣ������O�=%^�Lxݴ�G	��\�J� "�%`�M�	���P?��eHY�����aD>�pqN��!�kΔ ��'@��l�z�9W˙ֲ�#����}����A��ـ��qՇ� ��4��u"l�8q��X(W6����>b����s�4;TXYY��@�,}�h8p�|skj��?�s����g�5T{�*��AM�g.	{�����Fс��,<p��Ӛ��v�N�-���iW���JP\<��'1�C\��<�bZ���S�<�ZgT`��k�8�oٝjZok�G@F��?�
/�m	$��[^� ��9��A�ߏw�2�}k�x���X���j&�H��MV66�����u�w�S�{�J�P���:�������w_�z�`��� ,�9���H���J��_��_�0�q)��x�jd=��o"���ưѱ�(0Yԙj��vpPKb6�����1n��ADS׍Y��6�����#�sD�
��F��]CFN�da5 �#��thܵ�_�"2v��w� g�eP^Y�Ժg������n��`�=\���S��y���,{�\�3�]�4�#ymߐ|�!qV�7A��͑}CT�# Q���޺��|뿻��J��N�b�u_*�,LV	������}M����i�]�F<��c+�e�����s��g��J��$��Լ������4�5t�_.�B�O���.�I���������x髍䠒){�����:pZ@r�� 8fr��FJ>�������:;�/��M�������\����/�������vH��-�*�'��<N��M��FGs}Ϧt���ٗ����K�2�-�f3O�A>()�>h���2�;��4Y��{v	�;wA�i�q���{"�d+i<eN(l^?��ZRO�pr��I��w��"��虝�^�|��c�M��ӆ�L�d�zϺ�=NH�Kt���[ ��`j��WɴzgA�)UQJgq���/D����F|)H�I��t��[M�z�o�x%*X�н]���������"#P�W�;yFK�	�s�Dܒt� W�l�ʒ�J�IWD�~Y�F
pG+H5`��0C�К�,}�=��o,Ƽ�vB��z��y�Y��ڗq�%ڼ
U9��^>�Q��t�@�71�R�m��Q��;���ވN�q���k�3e��U���n�ƭ�0�*��N��ҒQ�E�	�a ���.�x��ݨ�F��ۦ[�I��RZwX�Wm㢙�O$�lW��A��}ccƸW�X��#�5���s�mL���K���r�9��i�V��(>�U9�tŦ�b���-A#������@M�'p |m�5��0����ͅ,��O�i��ưz�����	�4�F"����w���&Ye���f���l��+'+j��\��{�nk��z���捾ۋ��x����s��)<Z�r{�<�*^�C��Y����6u��}pfV�꿗�˭��ŋe��w����|�Q�wr�?M�ټ���3�2���=5\�$�ۣ�_(�9���R�:ce��y6�bw����`��;�吂^�`����&���iUk�`FQ�A'/�\�XK��b'��r��3���Ԗ�6�L�m$�����8v��M1ց$�E���r��(�{��c�^�H�qz���mi�|h,%,�ҏ�c�y�>h]��YS!��nC��_ �$��4.~$�&��:����\T�c�#W}���p����x\����U�gkk��^J�X-/?0�{&�g�^�nnO�Z)���)��_S��$dX�R'B����Ҿ�"��A��o�%��@@7����+�y�z�A�b�����j?�>��g)�K���a��!hy�)qsR\��H?��B�%��2����������-�O+��y��l��B'b�)����6�V#��R�&Co͑L���E���VG=]�D���Rm\X�^��ヮB��q�n[Y�z֙?aa��� �����$	��cZ�ϖ �;�oLN��#8�ް��#��$�c���iٮ�D֯������a/����I�F�m�\���{>�Tɼ���v2��=�4G�/m�D\�'&6v�V��Y����ƅˉ�ηusk~(6e���&�Gq�
�j��j�P�mOxRd���S�-s!��{mw���֠��h�	�&��R�Ȩ��J�B�
c ��F�Fu[mpJ�}��c��t����G���]����Ak+�9b��0����u�:�u��O�~:�F��P�6��8X�k/��/3Z� ��/�A�X����QN���,�ע��F�)a,gLҜ͋m�eNMQ֎�{6-8��4~	�I)�����ugk=	7�����~B��Z+.---Z@`Nf���ի'8\\e��:9���R}=>i$�:թ�N�U��;�u���T=N(�|��j�G���ԋvaQ�$���$���Q�U#a�&�5��g�U?��R�y�����I��1�l
���`𜓠�Y��:������}���Sl�d!�"�j%��>m�a�����컴�j��Q�W&�O���OX�U5؉�?,��N��r��~�������=?��Â�Ijj�(a�u�	�tkݾ���r���q�i��<K��C��}<Z�%{T/���]Y��R�@������S���]��R9, �	.懔Zꝭ��k������
�Ժ�/t[���7y��ҋE�R�,����w�kZ�椌����j}0���0:z�,Rd��[)KU76BGNqFùd�X�N�P�D>6���iX�����w��YI�'��3/���gTt���Zz��	���@�'��;AH�����\J|4��E���ke$,��8҇=Z_y$=󮤆L:YV�v�~)��9KM*�x������������\�g�
�Yd��_֨HE�cL7�1\Dd����3�Ϸ�?h�j8�iׯh{���,��MW���ò<����\jͣ��R�Y�Q:df篇�_�c.���mȝ�#lW���X��?'���ko��L�+�qzݼ�y0��`=�m5g�8M�Q�(�s�hx�?c+���2&�J!y�^O8�ޛ�	�0l��mT(WoZ_�~N����Y0�<���b�<fj7FC���>�����U����yo`bX�2ǫ$u��m��ܐI$�'��;��X>--�o�#g��L?k6V֜W������n��uttJu�����U�R�rq�k`���M����y�I���n���!����oc�(����|�H2yr��@X4U�_XP-��=Y���VD�qu�HØ���C����D���=��1�J�tۆ���cߡ���a+`!��O\�P�z����z��n����]�R��V�L���B3R�����.5[��b"��I�^m��++u�Yno�&�/rq�*t�Op0����/�<~���	�!��2����~�*q��8�����+��&o���B�����bd���j�)V�����f���S��4���ԏ��[@��ĉ�j���E�"|�UIqD�^���"�N��=�L�SY�~=���$t7t+]lح��ɋG�y�|d������8^H�MJN�]h�H[.���1�sϑ�Cp��o�yH�uWXǺf%>�B��K�^�rLp���skۜN
�E� ��GY�~d�PN���+Q���ҮI���ClD�7�bpC#�i��%�� K��E?�@��O��L�?�=��/N��?�w����7��g���]4B���ۏ�QR귕���R���Hp�8é/�]�X���8���ks����Z��s��X�<�
y� aw�	�	Ӓjy�_K횴@��A�ς����
�[k܁"�I��(ei���6�}�U���O1�X2��"�</�f �OP�w�L�zB�\�U�]�:ov���g���K<�+ǥ�N
�PH.�-w�N�x��-�ç��u웫>��N���}ϣTk�,i?������8�ʨ��%��%�!��wBp���݂}�;�/�}���wy�~�{�̽3�]5�]52¸��Ch�_!��V.%}���z]����M��rj�NC���%j+�4:����.^�J#�0!<~��=Q8o#�U��{��5=;���-%#��m]#��&Z�5; ���󇹷/���P�3%^=�;�1X��fS˽��Y���!�٨��r�3/�<{D�ԭ��w�"���6H�W�	�o�t��r�k���O�|���/s��e��x�P"��	"����!xg�.��O�&�F=;a�x
�d�{�7DѢܿG��"Rhk)#0��Up�r{�3����
��sZ�a����n�8���謨���q񽯣�j]P�@���-E�Є��O^��y,(��H�l�q��cHm�0�`R��^$�3�W�ʼ��Z��&����l2z��ۿ0��XXҟ��O�N}N��m�^/.��l]\0����rf�r>#×�o1�NZ|�,Ո� �MT��r�A�&Vak�,u	w{ݯ�����D��r�\B��,q⦫�u*O��t&ъ�R߁�� ����h�Rӕ��I{[�M��� �?��),8���|��bz��|����/h\p����qB�C/v/���%(�L���=��g럕	.���ľ1�eu��Ҳ�=b�%�D[H�ܼۻ4��ԿQh1E�o�B%y`�DCʇN|�7�Gן>��\�"��T�O��7���2����O�XZ>R��[���e�G:�x��~�c�c�� 7��M�yFY����=`!��3��J�Z�CD�0gru�E�kj3�픹� {�3��8�+�e峢��J��� ���x��w,sT�'q��I5��~��@�J�Ǟ��Rk��XXXP�	/�?`��4\���2Jmࡶ�'D�l-�?5hO��)V/�S2�u3�O�o�#h�8l�����zѮ��&)|��'t�*���r��ϐ:��-�j����ߓ��XYX��v�a��o��,nX%��'@.Ī��GX&��HE��v+o`�x y��:`�*�r�e���G�&j%��|
�_� �����w!�5��D4�p�8X�-)�$+�W��E��TY��zbzP"�H��;-h�{b��Val�g�qb{����-D�������+x����{�i~ޤGf�`j4):��7Ϧ�i��n�pX�w@=^ც	���v�w�v���&�0�5ˬN7�{r�$J��h��)��E��:ԇ���Z3Q�����;��kϫ)��8��CXhRM�7�R^�e9�7l5n!�Y��-���ѣRw;�b�xA#E�BػW������,��4+�ϔYvv-u6H��R���4��!��DA�E���[D�"QVe'4��@gM��w�),�`Y�����K��d��G�y�b|�&לfUL��T����iB�7Fꃈ�(�� ��?#緂f��"��Թ,$ޝ`���`�|h�ئ���/�O7ʩ��B�Q^�ș�C��i�_��W7c]���1?�A�����_���	(�r�к|�n��S���W�z=�V6�p�ЊJ������g"� 6%/�dFRa��/*~Q'z�J�?}f�_yw�i��/����R���7J'R{�lu�
��W�I}?088\��E&v�+��!��iX���o�z/?������T%+��\{�^re)�%�u�Z������	Ϥ�-)x��V轂����$���o��g��$z#ǈ��8��{�"��1�<���(��]7���#�o�x��]zo?Ţ�ayľys ?���#Y�7jlr��w���/�j)tߗD*ꔭY��C���"
����ơS�S8�Dj�n<.՚Tw�`�>��'s�ި���V��z{��cgc��S?����������Lfo�q6�~/ =����$!q,~�Gj)����W,��_w�B��_ۺ��]���D+㬲��U�f#1ݤ��,L9Rي����׺\��S:��j�x����ۯ�E�.��lP�Ki�L�<S5t��*�������9�������(�E�X��:�F}��{h�47at-|7��\+=�If���>��	H����tA�1�C{<i�[MUO�rO?��q����[��m����.\��{��t�)�>`i7pkkg��]�~�R��^��s��lP;�9pU9�/���t}t��4q�x�e��/��6~�L�#WE���;�4����'0��ԝ�L��x�7ʙ(��7_,�rM�$���H�>�^�f}"�M5A"ke ��Yt�B���b�v	�Ny�Jؿt⿡���1�+YǏ�Ȟ�d���k����j%��J�l��2�MɵQ?����Gzx��)��21�L�T� ���MO�+�b����.��n��+L۸q �!�YHqk�h��j���!J�D�L㳒����_��
�9����>�q�b�!�(��7uE?s%��G-��(
o{����j"g�v���7��c, $H�d]Ҋaw秽�~���ȧ��G�y���������=�p��~�z��sDM�T~�4�L�ϝ����a$���i^7�`���\oP�{�<�cd[E�A���.�d��X�:�Z�L��葑��p��D �V��k�/�������WQQu����s���3��":��uí��?������o�������fՁ.Z��~�˚���lQ���+��$�=����v���]_=��]��Q�ߣ��u��y�ʻ%�@������
-1,?Ϲ�'q eP"��a��CR��xN����.:�N��๦�3�����g	�v��këa9�	�w�jI�Ά��E3�vk�R3r�ɚW��v6-��eD�J����g!�}tw���5�s�[|;�۔gl[�1!��f�}�>]����`�'OXu�t��m%��Z#g(T����^Qk0�l���4��(�,��:ŵ��4�2�EFU���B)Y�˰ ��<���+9���4{��ˌ����������A.���$���VfԎ��d�*hlU눯3'ۙ�j���U�eߓ��N'$��R��.��)O�G����C�Ц��.���uukgs��F4E�W�F4������2_[�,ULX��%�Y��J �(��j�Ҫm1gY0d��)9s~\795K�����~����Y	��J�#Y*�_�ڭf���<�W?�$
�#�״��ҹ_@��x]���#?*^���U�{�@R�5N�籓���Y��	aA���}�qJ#�胋hhŷ������JV�s�$��%�@ ���Y��~�#����7�>������j����^��ۀ���^�л�w"u�~��QÑk[��[�VEe���:�(�6`��a6���-�.���z���l����+sN�N�#�+�/����8֯��f��3���:�M��6���c�����e;6vv~Ո3�������wù"W���g+��NG34�|CϷ���U A���r�t�i����n���r���Bm:���vf>���9=���d,z������;ɭ�{��i��,�����&����_��u�m�=)��OL�^������-�-�%�zFz�ς$P�d-N��4���~�4r�=��<���1��E��k�[	g�fo�B���>�45͠+�	��W�3XVo˒�,��Ǧ�k�e���':y��e�4z3��'���a�n߾(y��>�}�)F��c���\ .�/PF�t��^�WX�(� �8K����̢���@�-�$�$E���Coɧ��j�ώ('5&�3����a\N%���SbL$������G ��b8rO�E�J8��B���	\�U�0�R��|�E/�c<,�A~^�*?}l;���-M�����꤃����z"c��P	w*]�a��tAM �����T�<񔺓����τ�.��"X���k���l�o�,�ն��~)l�U���(U�d�������K�#fW5C9�&��}v��� �HqI��߁�e��|n��I�����%�/��q�E�v��3!%�;�
o3��z�^���o�n���**�,Uzn.�)������h���m�����5zѺ���cys���pP������7dS�l>��y�l���/�u��Qo��b�u�C9Wpt�l��`}	dK��q�uxn&t?�i�٘1,�^��\%x.:���(mViq���{�a���J�5��ꃊ�%׻��e�AF;נM�x���YFV����]��� k�5*J��j6[��]aT�����x�9 �Ơ��I�O��g��xxZa
��]8�L'��t9�`�>��~J�C�^�ی��w�p0?��}$����@�d����̌�#=���;�U�~�ro��?�(_8��lc��������Y�w�Ã��e�P�nY�e����
�1�ǌ��2�	!(z����3"b��!�r�/k��V�l	Xu���qn�o�GCm�i�(y�yt]y��k*��j�
�i�()��q�~(;��ȴ���˱AR�#?�͌���7Hy$N�%�O���z�ԕ�#��m�O�6P9w�;���prP+�F9W��5����)��YK�?�R���+a:�߄b���O��;׹ Չh^�Q�����A��W����t=þ��s��q-C`�Zު�I��*Sv��h��r.P�@�]�S�9�hm*�5���N���tO}<N�|l�y�Tu���RX9�&��iH�-�V���7<^����A{�'�.�Q�]�V��{�\���bb�K&�t;A�b�@�!_��e��)z�x�%>#�� �/`[��#���y���q�s�U�cdȩ"?�<LIz�T�Wwc
e�^���r}�~�N�nn)$�	�F~�ݝ {�����Ѝ�{s����F��L��{�w^�D�)*:��'xTe�g����޻�#Ν\Sk- ���Z�oH�-�J4�J1O����Xݒ��Gɘ�g�>g��A�r�E�G�)U���>�!ݐO!�cR����?��Ӎ
4���8�����c�]0k;=����d�=5��46����d�A�7����{�S�!��O� �������,V�0Q�!d������D����5�"A�����`�V2��Z��p�c�q�}��7��pU�"�_��J����ܼ�`�+^*��[Q��̚���rV�2�LZ�T��g���`���,�L/����_�T�vb�g�3bA��D��_�5���cˁ�0����`	4ҟ�,��Z����V��������7������/��&��S�4&S=�K�^�R�T�j�E��ݯm���3z�r�r#@Ǖ)�H��ɭ]_�;S�Ol,�;F���|��OS�ĝ?��$�b�MLG��αi�}od���R�G?�6�x{�%ؠgO��W)�d�y���8O�4z������bH0(,��bx���S�$|5�X9Pkެ� $������	��FR�K%Z:���,X�L��	� 6�=���;���S�u,��"i�uVɵ� ?�~��K���2�/ xC�:������Ҳ�(Ӽ�{�{�R�����sl84�������[A�7=��H7]R� �x8��](9��t�ٔ
�l�{�1�
��_Y�99%u������߷	G��k�HiU���I�n.Z��[�`�׵�[�t��
҇��}У+V��m�q��^cf1��vH��'��5"�?[�|���q{�G��1���fi��=0�Z,:SN���?�y��p�b�%�;>"߿G����,�-doŨ����jYjv�]ou�{���D��"�:��܏X�ؾ
����T�>�u��c�,�5�z"�xAi���ѿצ�O�M��r ~��m/ (+b�!��^�fQ�3)����J��	�՚4��!G���e�}������(�� �僢�7_ܐ6�h�,���s,!��2�St�� u�/VR�h�9�ٞu�Ev��[.��s��3˸z�E�� ��k��5�s"h}�@*앝a�j�R�j����5z@Q�S�%�\9�4���� �;��w��8�L=<I����I)C-����O�_��Ilus֣���P�=�x7<9�M1�����h�H�����q�]�
�����C���I���7�8ͻ������xb�\z��n���9Q>�׭<p�	/��q]�'��R���N�rh�xÝ�2�o8�[�N���y?/���2h'�M'�̘(���ndfay7wx�Sq,�0��~Y7L����ظ�����`�~m�XM�X����iNA�;���~���R� ��魩����6�)�ӷ돉	T{���( �����R�0$c9=!�K����</�Xg��E�h�
����k�&
�����~`�<�L��70�uU;��v�ۨ�ј�CB4/�5�}�'�k	� ==��C\�s��szf�<l�W���+�(t�<ϡ��mR��������-��eq�THD�u~��Fq�b���u��Qu�_��30�kID�<	�ߋ�)��$��'���E	�8LQ!?xK,�w� ������?�s��# �9���΂`/��Z�&^,���I���\vS���ran���U�]�yY��]�.��LP1)qZ�0��M盒�]���w�C�%���ܢ��N���i���D�iZ���F���7�KR��;�H�]}���}Wmdm���ڡd>��߬J����C�gvO���ǌ��fv��eH���O�gNܴ�{��3s�o8@Qer�Q��������c�(�OD�x4��ʬ����4�e�� ���L�od�AP���y�?33��	Ys(��. u0i��sѦ������J�z�^�ql|�����-}���hV&Z��چ�}k�jV�܋4ڼ�v>_xB��v�n�M�$�־u��q��5���M(��#��	F*���ߍ���lg�_��z�S��!�ˏ�V��a�PPVYYƚ�H���	4����ׁ۷)ݾ5S�c��:�U�-lJB�lY�gjq:�����7�Ԫf��,K��r��q�
8�-�wo>�P`ff=o�|I��<��0�OaCFD���F�@'�E�<�j��0w�4�^⋲�lNŢ�z�7,76@8�T�8@�888W�r0ͧ�c��,� g�	�̡�}5ZT}���U�6XP�eD��1�L"@A����C~����)���?���s�|V�(�<\\\�L�������Gp/5�dR����v���o�h�a�斂$g���6-֑N-��,��o��W��6���apr��vNM���Y�t�Ό���3a6^��@5�-�j�f�1�j�c]x^7��=�����Y�h�[o5��s�J>8���#D�F$˒�*�!*��	a�*-�9�#g167����I6o�&�lmǃ��=S�T��LM��KR��frtV��f�:�T'����-�;ή;TRa�0މSwKĮB:U[�SO�o�Ͼۓ�����9�~��	ӗy&�_'�����wzEn��z�X_���4���p����R�'�J�?�� �p�r),Ϝ�Y��z�PN�G�<;��]n�g�K���7^�|~�����C@��R��JF%�ݰZ��,B�S����|:����_b���q��>P���ڍe�5d~� ��94�x#����ڕ�i��P�� nIZ����~�X�`gQ�Lh��{0ٽb|�?X���Okvnm�U��"�qx����=�Cb�P�!�����j"oE�~%�ί.*�O�M�ʤ��<����%�Fe�상�0��id����"r;0}��^���s9�$~�N������zq-*-�j���ȳ�ʖpت����X�j���aӁCQ3���֙��H���������֑i�@�a�b�ecQ�8�]3��i���ͻ��j=M�	a�}����2���|�]�Q�Fa�1� de��m/x�W�u14I+)ʳ��3��0s��:hx�i����%
;=�<h���{ܵD��" 4� 'k�s�k�B�M�5�#&Hy���3��'I��P)�-2�����3�O08�Խ�Z�t
��a����D�J��Ҏ�h�$�	�XAg�O�Vt�N�y]�M�������F��0�/5>X68�΄����p��<!�:�Y"*�"�}(5��o��m�8�C�C����h�����V���;O^��m�����0o���ͻ�A�d�k�ߔ[s#����A�/���U���%v��^�)�ѤZ�%l,��>�ê#��wy�+-c��(z(3cx��|i˓ĶH��}�*�������`�[f!�Ս��i�L�*��-%ϓ����-{I�����e���O����� ��_��k-(b�n�K(���ͩ�3ˣ+O�-�t�4@g1N1��n��L�'�S��;����Gg�r{{�rՒ3��1f �sŏ�i��F?ss
�(�C���yG�^�&9�ڲmY��?G�6�V%�e�V�����x�X���^ �k���2+\���޷U.@e��ű�O�`-"��rA�뤡RN�A�'�K͍���)��r�� \�;���H�˼���z�ne� V��l=��I��l��{�����]PW����_���a#x���G���[[bȡg���T�ұ"}U��Z�MȒ� �4,<�4X��H:�.RU� �9Rr�OI�(� h&�/J��x��y�����|̀�k��K0�� t+�?�0��\�|�6�����h�j�2�_���bM��	/j���rX�#MÎ!�,��bMG��G�6�4ct���4��q���+�-�F)�~*����lI!�R]Dp�D��)�����s��@��u��}��
��a�~`���8�VM�J0��ʐ&����v�d�N[��4�Bc���l &b���z�����.���"@��/��/����f& �o�_N���A42��.�A��j��jYq��:�D����޺�[Z�CZ�� 7
�+��Z�E�n[���x�&ۼ��L�5�v��P����e��rs� ��q����-s�c[�j���~�5�8�`%1'���O�u<�_n�q�Pڽ�*��V��:��^#c�~�k��`��km0sE���8�JS߯�,��;u|)j�A�6ai7@)[~�0��`���a�M�� �� ���NE6r��*����7�b���ԝ+�������]Ym3�_��D�zܮ��,������J����c��c��pл��0�����6�hz�g�l}@lV)T��Z5q���,����t��xڣK_�LJ��/8;r �t���R�*��N[������@��ڀ�n��;}�(�'`�hn�1$��M�[�gi�m������I��H��	w<����gXZ��S?n���xgÖ��7"����0]+#u�Kuq2�UIX���QqB��:iŹ������;����LkrT�䬹�+���1�m�&'�W/�oB�Wj�=~��
��
�"�m_��ٰ�-C|L�����n~��,�@\�/���M���
c��ZIE�l1c�rn�}�0��m��ɳ���8�՟�o�Lڶ��t~V���v�(�f��st`�{��U�l�U��&�k}�d@ȁ~<��91D��u���� m��639^����8q���lf��@�"�q�<Z�*�*R������T�vam�$ �ȧ3(/N�1z�|��n����I����x|.�`�Z|�K		�]cN-�d��b�H|�������f�ȿ)����ְ�~����ߕ�4�<���C�.:͂Gue�j���Qu�r?�b4�WKV�P)|l�~���:��i������<�SDi˽�ͦ3�x�L1�0�H9��mO?�>��7����9�~z"�RP�����+�G��]o�xU�t�ôk�lu=�8�]���"�O�L8�!W�wk0H�|�F�d[���RI��dJ���+2�}GA��tN�U6��?��w��"����08nQ�\���<ʳ�1��"	�Ӓ�z�.\
G��@���os�9���z����00��.���ס���<��`���*�z�.H����IIm�M}��c�&s�Ǘ�]`�"��v� ����-�#2"���\���<ʌh���k�G��~J�>A��:��3���}��4���H��[����4MMK-�[<tׇ5h�5��}Ø��d4�d�F0�����U:�O��P�MT�D4�����i=R
}وx���h�٣�>+���e���mS�<��������D-�KA�ְ!a���c�2_�{�K��pGV�cN�7K�e�ᥓ\7ݓp���R�F��֯��e<�K|DJ��YT8qb��lM���~��t��O�F;�2V�}M*JI�!y�&��&�1H�G9�Ƈ���
�1W�t�|~���p��}_\r��)�]|�3�B�|�=O;B9���ʧ)Q$�?�##]_�*�q���D�fG��`�z��;��JY��Č�x�/dv�A�~2�@�r��J5��k�V�Ɩ]���n^���!$9�1�[D�2�C��)�9��t8���9bk���k��Z�9/���mL-�9Iu��{A=gG�yF�x�_�P��8F��~J��<V�����$2��w!;v�p�l��HS���#�
���
C��ضlϢ���1Rr��3e���[���(����q��X����mL�s@t'���z����Z�!�y��7��&ݝ�1���σ�Ϙ�%!G��+%jP���;����N������f^t�%~��P�M0�{��6
	��9�z"��O��
��џh���8+SL-� r�`��t`8o8D���H��x1q�������n���N��YٲH���nlS���f9{*����.:�i�ZĒ��s`��c�]s̀N+��Q�OM�74V��ڭ� �Ȟw��rm�� �QT��o�W���}�3N��\�O��4��g?���:�c$JVa)��LNgh�Oז7ڭ&wF���a��6�Ջ\�����������~x�3�b'2�>cf�9r�A�X����hY(��݃��5�H5�=T����j�N �=8��2�`�Vo5�\?@�MZvH7�?����0��d+?��2�%�Y���z������wn>���߱�CW"�Y�di�p�X4�V;S0_�TTWy-�ڄ�T���e��CI�&	��$R��}����leI!�I���,�����Wޝ=�6 ��*Sk�y�4,��P!���#В��b�#�։t��>U�J����7X���
)i��~�(*^�a4�MU	�Ô�GD=+��S�Z������a��WC�Gn��nu��o��ن62Z����~�+z5,�+"F'"�wېu����!�g����>@��- ���+����:�|�O�p���f�"��I��-�6�m<}�U%ǖ=B�I���~��cC̳.x��7p-^B�,�k�f�7�8�!m��ON\ȷ~:����"+�7R��C� h?��`�卞���l�XZ�/,���b��5���UU���Zz��.�j��G��\��oD�^ݲ�X������������^3tC���(��L�uj����+�+n��o����>����߀�6���	�h�֑��V�^ �QC:k��"x�,�S�W�a��O�6�NZ�h���'�U�@���J��寈�弾�D���x���Vjpmh��s����J&PQ��ΰ��Tʮ�M�c�TDF/HJ2P>�eN��(گJ�S<�7.�<�>�2U��(�8�8y�FQY���e(teai�|6���ήV2�f�´�A;*����V�z:��T�(�HG��[L�� ��?��EEa���{�0�dE��_��p�F\�D�%	��6b�腂[�z�ԑ�����
��.Rwt���������>���}�>&v�m�W*����|��b�t^ר�|[$rH\�?s&Z�{|<ь�E���w�)�x�|Tc�ׂ�|�QI�>�#�%���+�X��]�h��Z������tOb��O0�͏������k��D%��X��~���e���R@-1{�_W�-(�e O%��G�r�q}6	g�2���;�8v�Y��i����lJk�3A[����zߓۗ��>�N=���Y��Z��_�*Y@��⚦��߾o�w��T��)!�οtd�2���V��n�BO�5�t�Sn˫����nW#XD>{nN�#�����)��l
���iϣ3�"���#$�vY1�$��E,ХŌ�������>�a�̘,�#X��X�U��kR�Mv���,���k4$!C����wm��OӶ�~�H4���>��%N ;�J�|��6�gr�QM*��s�YD�@�Nv�W�l��M�3�z�B�}g/c�l�`�Bt�C8��$@�g�*]/�j1�����r��Y�9�Ͻ4NI���K�I0��H��Gĉ��f����?�vbÞ�������/N��}�R�_VU�JSDPʷd- �!���sK]�Hh������P�5%Q���m�G	_Z�C*�10{��Y║�!~!$\Kf�dK�)F^���uw��j�0|��)������� ���*s�$b�u��}��Q%�%�yX��}4 &�%��y/��.3�����ϭ2���O�N�X�h%��������fA	@G�k^�t�1Y���������f�A�J]�:����g�7�#o�����#�#tڴpz���^ÿJ2�s�l�z<���N�Gb�G����Й��y1G��-�?c�4R�K@n�Ώ�\��1`'�:He�fd���<v�8-�(�(2]O�2�K2�<c�1P��m�!��1D��Zo�f���L�v�#iU�0��	B3�hS&�����Xsz\�˦��;P���̏��M�lB+-2a��ڛ�s
Zq^�l��H�!�:7���A�$ݫ��$�c�"���ax֏ݏcF�̵�f%��#��1"u�m�y�fIZrr�����Ӷ`�l@�Z5e����q*K���{u��^�"��2���FX`�ch]��+JuA��W@��vĐ�
<�G��g�-L����M�K#�[����o~c��R"��*�� ��>����&�)���72\�z���S�Rϡ���.�r'�/�X��Ҙ?��WK�^��Whv��:�A��5�<��ؓ[�,��-9�`G4��*o�G�6���Q�`�ܷ݀��\]��d>� <�2#6��jħ��e��2��g�G�c-�-0�2�7��UAo����Oƈ9��r!��R�>��9�ru��۞�f���%.Й��8������J鏛�4ձ��:n�2b��1����%�f��ZT�� w=;D���k m��Ҕ���7�I��ǅRʋ���g��K�k$<�����he9�J"
��ݲ�2K°��l�mz�ř�P�����Q&ru�՛=-�M%�A�F���I�p�����������cq��hV�Y����I<�,۵���}t�ο��Eȕ�=���������dp�G$���[oa��c^�������-�����(��kp-����܀��ʂ�gr�`Ǽd	~�Jr&��c�j��4��d��)�G�A������I�v�EL\��M�����r�aE ���!T֋�/qj���m9����%��"��:�羹lhS:M���G����G�y����	�p���fGh�k��,�Ė�C7t�9�;���5|����i�=[�.�m����w�,�<W��i	��^�V�ؙ�V̗"w�Џs;7����k��]��-���&2��ήa/pH�%}Zh��U-r�Y�� 2N�ū�ab���!����
	��h����Axeb�efeݜ�ކ�9�m�;�_;����_����7|�^�h�֘ �i�;Oq�L� �M?i�`0�G}��dv�o��sO���ӭď�}fos�����Bf���f�W�.7�!]�^���w�
�m��T7;�!�-Gq[Z"䜝��uJ[��\3x�F>c�H�#�
Q�Re~��c0-���_j�䦓 �4c%q��v��+:���)�+���e�g�+Dd
6���pn���StU��h����f����S��b�@K�*M���:����	g|qd3dlWl���d�'�(�!��0Q��G��u�y�\C1:� ]DA��������2}h}���Ǡj�D$34 ���O�j��}i�-(�/�]{��^�
���s�ˀ#�Sσ\�A�^�m���?6���bt\}M��F�x�����*���\��:S�ˊ.)�V�'��^I�#��'~�/�(�S�X^C���Z��`���W�� �V�����E��W�&�.����!�w9Y/W�����T�����H�@�zr�3YK��5=XV��]��h��4jܢ9���E��9B��a׋���"n�|��(���' ��e��t	��J3�)�n緃���sܜV���]8RÎ�K
�B���]����[=b旫_�1�g<�q�9l9#�����&R#�9j��/�Zߧ6��i�I�}���;r?�&��/�l�I�J�?�����Ɓ|^�Z�E����8����Ov����Ι���cdu(��n������	�i����=S�#O��`oyͽ�?���_������]�Ӧ����h��4�;:o?=�	�b��n���=��"�e���d%���H�ﾴ���i�pp�uF�&EGY;C�R�M�gH�e�X�	��
(I��}W�1<O~X"T��;ܽTr���
CT�B�m��>���ӣ�C�F���+H ����K��bt��VCV����9��YY�d��B��a�,�Ϟ�>Z�f��ཾחb�v�-��nurl���b����v��~XA�&A�Ǻq^��/<eƣ�š���4p��n�@: ����b��YyY�(��q��Ej�m^=�524���8��kfk��ۉ���B�DM�4�j�ÔV�����=y��>T��l�e�|%��}�����-��ѭ�_�ۍ�2���BBz��&]O�䩰�R�++�ׇ��%�ɵ6 3GR�y"=w��/;��+vEw8�4-��<��`�݃|X��z��~'T�M�����s��f��阇�������찬�q"A?�"�[D�H����Ά����4�~e�{�A�x�&��%N(���|����f{�X�Dٕ�}��׷�RmHҔ:�^��W�@H3\�Ɗ"'q�֨���(�*r+4�w�w�K&������xPnm����������Ђo��v�����
��C�zAa��yߋ��J�ؠ6Ӹ�@LN�0�����~���2c��
���[��a���d=�����y�cX��ل�{�A`��vG��M������o88�q#���vw�S]�Wg�a�I�F���y%J��+/����,�)%����ү����j�o����cX��08:'Ѽl�ׄN����	�r{%>�Ȇ
���OH���}���([d���T]���8�{�6o�æ�}�8��#�4W&zH����U���~�?��)�6�s��k~�zgاT��d�˭V�

��_��fl�j:�S��eJ�v}4,ZC�s�����"��E��@��S����΅I�.d�)�i0���9���\"��D��'�����Ynۃ�,�ARF��[��;_w��;�bl0Z5������z��G�.���V�:��ŋ3KӦE�r�(��q&�����γc
R� 3�g�`���s�ʢ8Ml�qi�$��k��r�:�}=��������8��;l��ڦ�� 9���^	���l5�"�/����~=����qT�a�c�5QW�0'����}��i&��Mp���H��:������0�b��Jqw5�p�ӷ�Aɐ�@ɑ�N�А���]�Z�AŤ8���mTaH�j�HiфZ\�����пE�vf�{��R�W'� ���G�s�)�qz���1/�4�{�mD�d����zD��6m�Y��
4��n�ӢA�Ļ3��(��cƄ~�SE�ϤK"��<!�2܁Ȟ��q@���P�x�n��,-8��yo.�%�������0U�'��4x���x*ԩ�cz�3�mlӯݘ�*~�a���4~��
��V{�#a���8-9���O�J!,'�H�
�����h��n�>��$]�G]�R0�xl�ѕ��g�'f��&��8%�_L��땔Q��,ژաQ}���Í���7��U�l�Sط��п�B�+P��3h���T`
v�1���N�{N kWQ�:>J����>�?��	w$�n�#�J��CP�|��]�Ga\@�Y�hR�"H��"�x?�z�e�GP��t���U����+uYS�v:(W��w
����D{�Gj��}$��{E��o�y�/���U�k�xN鼎��N��P�ˤ��m�x�|���X�Ģ�oHͤ�G�nD^�G���4�sޖӊM"30���F"/�v����s�F�m�qC�=�S�6���C��s����3<���S�ZnhG0H��@=��%%	Ð,�زu+�.^`j�ޯ���W���EQN^�a��||? �2�$��=<!r�,�Jn�?��Xa�s��Z�xүڼ����g�˵����v�fl�5b��zpE ���o]�(�sq�����R���D*E^df�̙�3��ӏ�����O�L��:/d3W"`����S�Fkd�L����D ��V������j�P�ٺ��=a�l@�0�`0��Pl0���-G���Aӽf\Niಿ����	!Hӄ��8�w� .\ �c�6�}[tށ9h���+_�A�|�N�_��|Jq	�yc8t�ۦ�8s�8��'�u)�%��K�/p��9f�gغe+� "K��� �`&s�QQ�G!ښ�v�z>�:���h��� `��M�S���èQ����e����)�j�x�f � ���)*��?�9�
ewn�z8vM�(&��{�$��<bQ_ӛ[���/��ן��J�.׉kU:F�E>�;������Nd%�z>VJ�XO�Z
Z�6�R�ŹK���;�&�Fc�`�e)��u��aNt~����-�ˌ����>�v{ ������o�]��w����n�>Q�ig����~����X�N�R��ܜ��_��/�������U���F;�����=�\-$�}����a�I98����|�s�V��q�W[����ZI�Mܻ�$6�(�
�@��}\?��^/w19��ȭ���rd��:��Ye�7�������JIޙ��;K�k��H䶝9]���E�YJ�����UB]ZZ�t���֘��N]�=�]֢_5R�������[�x�9�ufv�Ço �2�ɲ,猺�ŭ7�wyg^��n�>���"}�<�n���v��ф !9pp?[w����7�K1���j4)��`-�.\ @�sf���c3�'$����B�8$�M�,\Ǉϵx��)oi,�
B#	� �i�(�v�!whl�4��dh��.J�!C�-C�;�u��s��ւr�m܀�X릿��<鶗a�b�����e���\�! B�I�v;t�m����ƚ���诵����r�,Ǟ~��WO��2A�e�ȧ',�2�g'���r�֛�ؾ��WdB�� �^�G(���8��������,-.���v��5a-J��7_P;
��1�)�(W��y�z����{y���sq�z��n�Hq���պP��`��0$���;H��"+�Ӥ�(bzf���%n�喵�����U���jQ.W��A����'���Hz�x��^���N �k�~36�ۏM��.�M��������Rhm���5C��,�lR8`jr����7j(�5 ��1�+ �4I�7/�Re�/�^����߮����VWW?��������&�`=�Ѭ�2�e����~��-[�����ZN�<A����<�4͵?�Poo��HA�O�V�cy�'8v�?�O�1�++L�̢3���۶m�ĩLl���(�ˋ�]��Ǵ���<��c'8��Q�2��q��*�T`,Y��?
�=�f�!\�^���X�u<��H|�\��*�-h9�]���Y!=��9�B�k��!z����ƚ\��I���v�t��ͧ���k��>ߏ�=�6���!�f�i|��B�@<!��J��0U�^Z�/|��ϽL�X&TD��L�hb��jl=��﹓��;1qH�fx�2=��X��}�'��)�~���,���*�.]��l`���l�$	�j��Lx�h���!���/I���<�GJA�f����+��a�;����z��e�]&���x���]w>� [J����Z�\�`������7�z˿_X\�HA�RkPRf�|�Gkw��>��ڲ	x7�=6�(~oN�,�u����)�sZm]�P��V�n�3�pX/Wp(@iѱX��2`2��+.t�c�)�\��6y�V�Y=Wܥ�z��p&����G).!�%��ϵ;miu^`g�R���:�M��Rz��yY�)����h�f�����ɂ�9����0���[n���r��1�I��v��x}���3��9�U�ܬ|Oa�����<��Ӽ������k��g���z��22�������{i6����跺Dʧ�hq�[/��)���uj���q2m�����4�T�$�f�)(E���^�ey���9�1�"Ȱ���vq�g$4�x�Ra34�`��lq�d�3�r-g�R� t���Qq����Ĺa0���V�Ä
i4q!���L�O,3�*1���ҽ��+�?ŋ�=E��fGm�Xx��Xߣ[	������s�}�P�:M�W��Ć=��B�	C�ߧ>>F�\����<������/,��v	����a���<�K���c�[-7��2�ƺk��N��e;ׁ��
�N���k���B��J�lX�:���t
@H��{A����v�.ޭ|;��3>6Ʈ�;x��xϽ������7�\fmSx�wE�𮟏�.��h��]��o�n�{l�wQ�0��(�_��aM� &���:�H��Y����׳�R)_�36֬g�@;/�qF2��Mv�6�̀י�,�H!�R���/,//���������s�18��1����/ֿZF��~����V�_���O�T�V�q�M7�����ӧ9{�,iΛ��+y}���#A ���VcSSS,,,p��I�}�Y>��عs���5&&'H��g4c[�I�e|f�=;vr��w#���E�n�&mv��1g����h�^m����	��� �xB9y8!�-���r����g��뀒 hO�ɜw���a]UI�T"�3<�1Zĳu�]��ͳ���+���{�e>pPB��� Ǆ�ʂ��6��`�Z��н>~����1/B�5Y:~��/��+�=I��%ҵ6*3�R����:3���޻oe�����Wid	�aC����St�<�crj�N��ɓ'�ַ����F�ݦ��:�cȲ�Lx��Q��x9^}����(:��|���
R�A��߸bW=bG|�A�ۉѵ/{�F������%�����0(���}��*�z�N���ZC���O��{v��$�
�x)�Q;U���������׈M��.�M��b8S����vYF��y�y��P���w�=_/Z�üN��X�,�����.T d�\�H�8��H��WJ��JHz�>��gI�ؓ'O~,��ejs-[h���tYX��������fl���:y��G}' oELNN2==�����\����yd:�Z��b���r����h�*Ug��������^�Lg�������;X[[���+FA8V!�C7�=9ξ}{��sg��\Ye�V�$���Z]�.αpi����6��kl��uF%��մ
}���|�ae�5�L
�#���c�}��t����X��<�!�Z숭k�=����q�W	�0a
O(���&V�A����](�U��]kग़���>����{�o>�g_8´*��	�0f|b��$©	?x/[n;Ly������D�SdRb��K����_��~�#/�첛����>��*$�Ͳ!g���i�	R��dkl�dhP��gm7�9����Fg��o�z�G���7�`-ښ\fN"=�J��������c?�c�~�W�/uӬ�OS���@F�\�f�n�f|;�	x�EQ:\m��=�-�ˮ��U��-��ZY�Rx�M��|
�S���� x�6*:KG ��x/��6�<�1�<���"���/���FQ����WYK�eHY��0|�syy��VWV�����u�|^��"�~�6��ux7~�N���R����$SS�<�������vR!J)��6q�̣�9�w8�
��($���R)�d)A��nu�u��_����ƛG��O�7޸#|J�*^��	��e���dzf�������ss`-�t:�Fk��_dqn�-��)�1"3H�,�6���S�p��I�	�t�jV�����۴:��b�d�+�d^�8����* /��]�d<���,u:�J��+�9�-6+,�w������k	�%Ԗ8����T�G��E�}�E^y�iN��Qb�)ը�1I�5ki��C����䎇���M��Nғ��N�q�|z&C��d&ejr�^���/���?ƅ�g����n�8��][Y��[���@6b��j�$�R���<�#Zg�a�$Ir���FJ��8���v�pvW��`W��f9Q)fbj��������&���y���!�ˆKyU�k1��q�c��������].�Qt�WZ�i\K���,�+���E�B?0�S�1���)䓙�* 8Y0��Z�(@��\���Q-�j������gT
g,���6�M����rUC��s�ϳ1E�\�A�1Uϓ ,R�����ӕ奇��/[�&�v`&��W'�`}�V�#\#o�9�����Az�;�!��>I��3C�LNL�s�.��<��N�'�/TCk��+�3����ͩf8�f��$��5H+�<�If�mᙧ��3�LN�r��Q�=W�/%��O\���cae�\�:5NP��ZH�}w/�������
���q���^DU�Gez�M�Ke*~H5��4��O����9'+0��"�+`d�<���H?ē��W=i��J�z�p^����Wۻ둤	Ab�/9�����M�&5�+��xB!�ZT"*�g���JD݄1��	�������G�d��Q*����Ee?@�!���o3}`������փ4Ki9b�צ�S���_*�d)BJ�R�'��,�_♧�⑯��o�3�[�	���h7p3�@C
<%ւ0�nw�GA��hS��������g���U�<������XdΡ/��Q��Ï3��:GE��r��0w�X��.ab�%� �T-3>>���%~�S?=w���e��[���s&��R��r��Ay
r���0D��b]H\�,��۩_�����;�\�כ�w3�w�}�`36ƨ���[\���}�㷽�<+,������䠹�BRh~
!s0�1Ԉ��eފ0y�m�\���I��0ʼ� ���������՛��"�$��¾�[��1�����=�4s�u���Z-Ν;7|\+�3�Nv)��`}�҂i]���l25=�����_�+_�~��&S��]�|���	��S�k�՘����s��X:s�����	R[��Oi�]��OLo���=�رqX��S�ȧ^�ray��Z�0�)z��&A�� ��O-�H@�����h���t��s�`DA��ǌF[��
=g�`���>AR(Y?Ay�#,�¯E���f�@0�xV�#�P�}M |d�!�]b��s'O��/�ZY��lQ��8�P)�!����j̎��o���=�؉���ud��W��-,/��yFkj�
J
�&���׾��~�׎�
�0V����Hz=F�r�
����*���|-�� U�8�R }�4�l��"�wΆy���kc0F�1I���,#.GL�ΰ�����{�ON�-d�,!�J��jM�&D�[鲇�����fl�[l����
)� ��<[���u>J!L1�Wd�$`ڣ���fy����
A�R杜]��R��Urx�V<��Ν;�{kkk1��	Y��q��
;��b��N����JB�i��{���LMN�j�X\\����6\���-��L^E_ ��@ �ŵ��b�@�	�X�̩ӧ8�{_�����O������w܆�$a-F�5/L�Y]\aj�Vn�����Q���kGI�Mt��L4�X��*��s�}�8�OO�e�v&��r��Ì�2S��I%�mFSJ:9��ٌ��@gh7k�)�$��@[Ků���2
2c\\�tfρ"�]��1HO �O�	P�A��%���-!�}��V0VCe�hT�1]��[^����nwx��y�N�aen�Z�]Z&Ra9&B���
�
}���ｓ��3DcU(��E��'�n���X]^fvzr�������G�3���.���v�I�X����)�#�^���4�\�h�*Rp�m.Q7������e���` ��cr��G��� ���Je'��j�K��/�v�m�"ӘV���N]D兓R95��4�flƷ���wQ�ws��º���:)l;��� T\V�6Li�yf[�U1м]���Կ5��l�Û�'����+��K�m8��!����,X/@+��0>�����j5t:�I5����q��j���W��
��e �Z���4�����ѣGI3g���.�x���{�C���g4��� ���r\������-�݄��cqn�?�O�O����I?���s��5&�fh��t�*c���p�0
9ա\.���Ð ֲ87Oky���Oq��	���Y�0��ePc"��$��W()�� �HI <<$�T��/]1��X�L� p4	$���M{{�s�J�3���@�$���Z���2���k��N�de�da�ƙ���S<��G8��Ѝ2��n�mӳ���Q��#�%����e�{>�a�{v�O�Ѱ)6�J��ﳲ����h5�L�י�t���O����7�řS'����z�n�E���{�()�-~��C��(�'�1'c�3%?xߌ�����ArU�,�F��HQ��,φc�u��mnTS�r[�4M���ĕ2�S��ǩ��q��E��۫���������ג$���r�~�a��|�R0�EP2��rJÕ9�n~������S6)���veY6��T�9���=��C#�5A�i�6�
I���ಉF��9�5��~�4M��`Hӌ$M0�૜{�eOz/�\eY��>sW4�~m��:��u�V*'6o���h���+�A�l6oz�G�����������K�˯���{]@v���۟1�ZE%n��F �|�M�Z|�#�c����c*��r��rI�,K�uC�����G�� i6x�OE4-�$a|b�Kˋ|�'~�_���p��辰��S>�N���JaL�Y�[ m��{�~Ho���W^�^b���N����W&�Pϧ�j!�"���ݾ��[��6�*G��2^)b��&(��kU�(b�� 3��RRk�+%�&���n����JW�T�3�=� ~>��'$V�^�e�H{��||��5i\Z�5�Lge��gΑ�6Y<{�j!���n*�J�D��<���J��Ϯ[3�g��8�z-��G�j����cmn��L`f�'���DJ���~�/}�K�]�H��!Ct�w�sJ�D�B��=�4�\�b�Vp�����j8ź��t)�0$�\Y��l��ts�o=�R1�>�����bQg_>pj��Rž�(BI�ߧ�i�V
�(d��]4�mZ�6������_��_�[c����J�$�4s����UJ\)�xR"�u�t��G��GZ�ь�w����������xw�&�}�&�}���Uf�uPj\����I���Ԥ�ӎ�Rg��c���b��
�Eq�0�:s�^�9.�^=�l-I'!C��+/���}�e�Dv:�[�ʍ��i�n �,8ʇd��}ki5���;��(������q�u���>Ug���T��E'[t�ŵ(*�2�v�S�~D��$�2�''�����=~�O�O���޻�^7���H�aSM�$�DC?%�������p�"���2g�������*��P�Clҧ�k�Z����
��	�z��d��S�ՈJ%T��a��:�+r@,�5h묄��'K�*T>� ��4[]X�R*! ����=��I�ˉ'�֖�Y:?G�l����Z�6l��$CfA1hk阌���r�]��u�^�X���t�4���}��F���F>c��JcR�����<���gx��7Y\\�V�P�T��ڴ�m�5�KetΛ-������ ^� %���}���kxv�]z�^>�.|���AN���Ɛ����}P� 
زm�z��^y���������N��ߗ��h4�|��ZK�R)��$t�]��k��h3x�.��	x7c3������G�벢�@HǏ�}߹be�Z��튀t���r`�	;�"ea��PyG]pX�,sJb�.ZA�\"C�w������7��ɓ�Z�8�(%s(9p��+\S(���{��'ȴ��LLN�!ǎ��sS��:p_*��u{@^�(E��M�i,.C)s����5�4U;@G�4�(���Yk6زu+�f�n�C�c�������/�~��K寰m��&̭�����!��kt�a,���wsמ-ܣ��&/>�-.;Kky�^��)�<�dʴ������E�,�
�Dq�\�|�r�����c����Ǐb|�'�D��',��A�ƒ���U�כ���d~*�V�����:]Ο=��yΜ:��y�*uJAH�ۣ��
YFُ�,�1�@$���(�ǘ�u���������쪯|�{�+��};��V���� �Ƙ�1��q�6��3�8`�y�3���i����x<`0�,�HRK(�Z��M��Ľ����u��� �Z�9��uoթ���ڿ�~k��ٱ��o�~
�Q��Dy�V�*7��D�\c��M�����u]:�6�˧��?�>��Z��6�J��1�՘,ϩ�B��n�G蕕��{R�������@�oI�� `jj%;�g�O�����bCU� �6]M���QV4*�*�^�����{+��I�n�'�Vĸ��a lt9����<�_�Tx��0��c�9�^�cEޑ*oQ�-n�:��:ϋ.i��r�$&Km5�*��4Ip�N�,�ȋJ��5�N�Z�R�k[��Z�8.Z�iF�d�{���MEi�����o��?�s� R�z�������u(���,�����d�x�W
A����s饗r��a�4eeu�J���,����טsC��jw�$�ͬ���q���ۺ}(�/�cj�y�E��f):�T� k\��D��=zY���?��x�w���n�)���M}+�0�J�`�ZZe[}�O	�K�Eh$Y�O֋8��~��:K�D�A�&�!ɒ������~l)�1�n�P��<�P��P�bzv�xY� օ!K"+I�Ϸ���N��JfHs�v��ۨ�j�<��0=5��yt����Y����x/�\w5�w"��A5[#�H'+��<Q���*s۶���r��j_|��|���{�������7�$I������N�!!z�*�i�^s+�5�0!�*$	�Tx�ግ������v�8����l�H�>�O��keMk����R�R�V�Ҕ�`@�)hLO�}�Nq�Js�����?�O�X\^�kzz� DQD�^�~��6YZd玝xc%*�G[
�Їy�?�M���>��Ȥ�;��dL�_V�Wh�M!㒅��\ӱ�H�g�f�r)�´֤yF���>�$%�͋�]����m�(z�Z���Fo�%�M"�e,��:��h�����������g��Zm��h4��{cP��B�� �H�v���T8�o^;�g:�q4�Q����/�K��`qq�S�N���i,��}�-4����0��<�]�����.B�0&y��;ci�y�]�0��%M�47D��
jS~����n�:.޻�f����*a�cX]lQgh�t���T��N���HZ'��9����Ӝ:~���N ���,���$Qߒ9�Ah+�ABߥR����ı�~T�U�$f��<�h@� ����ɐة�^�K�RAA�&VS�B��h�]���˫+���F���m���bj�N��މ
C��$�001������p]w8+��fjv�V����<��<����>��?�1:�K�A���k3�P��&����6���(��[�5��fyNV�\�~��Šw��d۶y���͛����q������G�|�Fg5t�]��q]��QDz�q����Z�?���<N�>���_��/��ʟp|/B�di1�3M���Q���Ӎ�k��Y�=�N�s�K>>����ܟ.�/�l(ol����O����M�40!�|Y�e'�c]�F�a�e����\�e���f�HxE�ɝ�Ut�<V\K=��[#�eek͎L�p[�[��ֹ%FaH�DQ$��ؿ�Ї>�_��UE��<��H���J����d	��dfYN�$���2??�`���8lJ;�-�����r�f�p�P���>�da�/6ܰ6�o�I^��Rv�ZB�����2�]u%���o�;����p�,g����=�g[(' �cz�6��I���R>����Q�HsV�,r��QV�.�m�t{�� i ��C���W,�5�;D��T+U��>���:��H�#MS�6�iJ�(G�8
�8HG!]�:��,M�T��f�jU��癚�ca�ND������.����~�!H�!�V��S(�2��m���?ÐN�C�:t�������Sw��)B��U��g�Fo ���KAx�l�q@�#�:�!3J�!�݊��LO#�&���}����ײѣ�u\r]���z�g����fiJx����A�#�s�cfzǷVdg���|š��������~Q)f�#��J@�:�A������s�:7�u�#�	��k�;��_i��H��@k=�",IoY!NejC�Y��4M�J�$˭D��|]�w��z�w�
�4��v�ި��}�{����_�/�f���Mk�^��(�RNPV�JI��>ә�CH)8u�4�v{��`��*֧�EQD��dEzۚ˄mN˵�q�)p������<Fx��lU_g 1#q�27���o%o|㛸���IS8��%M
��5�^�A�����d����PB�II��"q��'$Q����9u��V�#�%	F*���
�^�걍$zݞ%�B����X����p��'H��A2�|f�f�O50R��!n�{�L�L3�s������Kc4�L9$n@&���*���"Y�um�y��')�晪�I����E>���;��_�,������3L���A��"'-����cI[^=�X��͵�0�,-�F�k��V+�6�m��f�I���Q�O��p������)���r����=�++K TjUv�څ��vpd���~����s�_�i�WV���~��Wc�@K��a�۞	�`�'�I��_s(����z;�[Q�� ��ޕ��q~�YQ9-u�9c��6��
���˘S����"�1R#��i:��RR6_��_�K����$q�J�RNA�5�52;�0����m�l)�޲^��{�n*�
'O�`ii� 6}��)�N�a��T�,�ɋ���q����/�x����M����h�)�@J�69i�Әn�l����j������w���|�73��}�˵�^G\�W����B�
�HR��f�!�\�~�K�ip��Y��2S��ݍ#W-5ɒ�Uϥ�x���V}ߧ�]�����!)r�(JPʡZP�C�V��j�Bv_��Z�F*A�Bu���DQ��<�^�Џr�<��%5�d	�vO�c�������]�*y�y�����{>q��h��$IL�(G�0DI�T���i�Ζ��c�<m��uSa�c�k4/d9��F|��������V��g?�Q�X�Q9�3
W�&�4͆���Z�2�"�$E��nA��4%�2N�>e~�'~��/�󷫭�kU��zC���(�6�[�<Ak��8&�`�'�I�w�/+6l�%�US\��»�B$PC�AV$�Co���+I�4ސ<ϳ���VN�5��R��g9�I�UTcQM�� �wǈ�«sm�߇�c��QL�絏~�C���>��BX/`���b� @9�,������ua����;~z��^{-W^y%����������oT9zcu��=�t��}y�8��xp�X�I�n�%ߩ_Vm�ЖJJ���u�����O�; Ms��^��v+���5�y�F��gW�1E-&�)������V�gff�w�dq�+L�=�q�I3<�oIW'�9�¤���t�8���j5���l��چ�>Z	��C�&�؊������V���� N���K!�3�aH���z�tq��Y���g��'>����G��a~�,�N� ��y�`��U�0�ޯQ�_4����٦�¦�ؐ�r��!�Wh4c��qy@�[Έ��
��?� �2�r���&i�[��J$Y�r�P��WB�,EMy�Z�����,..�M�J)D\~ƃ  ��h@��Y�9����A�c�155��� >�%�]������~���6�qp}���)mR!����đb]u��0{��b�H݆��-$C���֘Tx'�jƤ�;�3C�1@*۬��h$r����S�PRa������5f���l
���@�T�K��Nk�z��=�y?�j����cjB�a2�(�۬B:���>ؾ};�F�(��]�D"�X/1J:�佘V�r�3l�'к����kV��kR0;5c+�i��)��k$����3w�;>�q~��~����r^������=��DQ���<+	PDkУ�V�k!d��L�u�Nr|'��y�3�^j�׭W��:[8�1L��`dJ=IR�4EH��}�BCZ����h��k� NQ����Ja�ĺ_xZ*41�Z!�^�Z�jg��˧>�1>�����?J���q�4#�]��&BhV����3�<���
�t�vN����ׅ��:*l�R� � %�fXX��6����+#Fɮ��J�����Y��86�7�p���*�q2$����>n!G1�m.-�Rɡ��Q��HOTJ�j��t:���[��������h�y�2����� �햅dC?}�	&x�bBx'��ƺ.f)���^�R�{!�V}�G�N1J� #tᙻ&#X��7�q����r�|�geu�����y�}����������(�7Q1�6{^aF�l��zCi¹U4�6��t������m�,����˩ݒ�~9a��ĵ��yΰ*��V)�(\�n�#q��^�HA���Y�G>�O��߿�������v^��T}�7��ݘ,Mi���Y�#�)�p���G8(!�u�4�m�J@�),�*>y�RQ���z����u�u�c����dQ�f�%��]8�&��<;pJSK֔���koFӨT<���r����{�}|����$��0�uϨ��%S�� �uJ�Z�z�iʠo	�̔%�Z���-�ѕ������B��ǲY��<ߜ�Ւ�1��[��\e� s�1y�6��hz��6ZJ�r��/gRR��J�ko8>�y�h��Q�XG�4����^�m��5��+Ͷ��n���Q�W9��bgr�ZR�]@I�1����N0�S�D�0���ܒ����͌MK��$I��YC]`�������v�IƫSVҠ�Z� ��C��I
�.��)�B�^m�>�n�����?��~ꡇھ�j=y�$g0�i�Ju�o���7݌Cy�Z��`��;��u�u�lt�e�:�c�^k�0%�%�4�eӞ}����>��Q�~RZ(�F�B�ϷQ���d�>�҄n�GP��}�v��u7q��������v�m���S�}���>ϙ�N!������D{m��z>�YJ��@��G�%8������&��W��"!	}���*�R�q̠�%�bΜ9ɣ=�]��$=�0�^�h!�U�8�	=���6�K*z��jH��E9
)@�Bu�y�����c�Im�M�%6~���������Y�Me���9M��˺�8 STq�ƭ��+�D(EP�	� ��a�%��q�ߣR��k�N.��
v���u�^;�+%L�N����G���~:��B�\F�%�aXAHA�Vg��y׻��J��g&����>n�d&�>=E4������3�r�.�S�-iЌ�w'��	&XÄ�N�U[�9��(6��4#��.,�֦G��s�r�>q[Mo�355�1�v�؛�6�v�G�0~�q]!R���*֕���ZOx׌��8F!��^Y���ɰK��<������}�{�[��ӧO��\pG��^��p���V*�4j6��uI(��� !�:��r
�u��9I���n��<r���2TiU4Ѝ�P��98�Td3��f�E��F��6YǰZ/��.����~������ZT��|��k�o窫�撋/�[naϞ=\pх4z�/�IN��`��dk1�I�EI�P�VG�U>��-m��E��r�T��A��tYY^���q���<�أ<��C,�=���ŵhْ0�b�d��b�0$�e"�}�Ћ�h�\wn�Z#ب=�]�f�d��`��q�R�vh������+��֮�r��X�a@�ף^��1�z�4K��_aX)�$	R*����ܱ����\���Zn��&���kR�Qw���5���E:ȇ?�!��x�QD4�H�{.�R�����K��y�-�5/���j�?����ٙ:�M6,gsV�^��cȲ5F��#��pa8�gP�1=��g��cK��41!�<L�_U�����	�,�r�){�^�KE�I�h\��z�i�r��`�u���Iӌ���Rΐ<�fE�둦�|X�ɲl��f��.+�X�h]������?�y�$	����f����(�]�Q))%ժ�|u�R#���8&)���ĳ�N,��Ð�kz���|��R�"�l��Kc�ȣ�w4Hcr�q����+b�ڻn;D�����]fE	BI;xQ�^�?L��]�^�˞={���K�_��W_��\p�f��S���:����W��H����5���q+'Ȳ��g��j�X<s�V�Ž��K���̙3��-��E��U����Lڲ������)���fx��^��>��m��ۙ�����nExK'vb��֝G��Z@�&�ܽ�3g���>�E�X��2�&I��o�k�╯���n{;w��q]��R8���rݷ�11�k6k�v��%�=�?�A>����C�k�Nffg9v�RX/�|ۿm��O�ԷEq��~i����7�s�]Sj��t6!��S�FgI��fH&�w�g0&�w��*|�	�S4�8J�a�ٴ��EC����F�<ːJ�s���������U�n
��E*�%%�UJ��*g���9���.?��3�N�Ӎ?�O�$���ǉ'���guu�j�� �Q�T���N?K���W]yW^u%�]w=�0djz�0�u{���p��iVVW8s��P��8���^��~�}��g~~�<��F'��I�� �lLr2���6'��^���n~K>7�]%��ƞK5Bx��V^I������r]I�tA�BV����^�bnn�Z�z�NV��j�a8����@̶�~���8���E}Μ=K��{�"`CA��$H����.��glY,+������5$VO�����f� J�'����tnOB+�幬Ԫ,7W�V*vVG��aLMM��[o��׽�u�r�-LO5�U�r?�%��a�h�X_�B08y�$�������p��qE\v�ӱ��o�������_��k�R��(�|���8�A�&���	�&Mk|MC�5�F���Xieoh���i��z��b�Y���T�����/���Р^H��#%���.-���~�����DQD�^�̙3�B���>�n�F������_�bn��Vn��Fk�T��c�y���qL�g�A� �VbaR	z���s��G9t�0ǎ�������?>O:��=w�1��M�Fk'���i�BJb6$}B�x��(f9Y��AT��>bvv8R�KI?�3i����,�3}� �ԓgf]j����毜f)i��m۶��|��:���.�Ч��Y��8�ܹ���9Q?�wd�觇�[�"ϋ͈�f�/��Y�L�I��~�����t�X]]e�������]����t�M��ʗ�y۶m+�4�S� P�Ն�kF �Q�|+G��W�e�0am׮]���o����~~��~�?��?��n��>sss�YZ��z�_^ߏ������;f�t�ۡ�k�a֎�4���<UL*�|Ua�
�
�x�WتoVh(K+��M!M5gϞ�^��ʘX��-����C=���K�3sx�G��6-�0�/��]��
�Et��G�v5�h�ʋפI�������P��f>u秖��w�x�ǆ7�J�B�ݦZ�r�M7񲗽�+����{/dn~)Jw��R5����+�;F�"PC��e��3|�S���c��9s�f���zz=<�]�\7^r�����(Z���VhT1�+�\װ4����Zk�Z�
>e4�y�9Pui֯�P�G?��
�_Y�����F�s��ژ4�L��Έ~����X�g�a)�Z[��r�:ۨ����sUxG�Ƭ��k��A�Z�Pz�1��fe$��g��r1LC���"�J6BIP�n�����J�����W^y�nc�v��˯��h�v��6����Be@i�E��l����޽�u��z�ڵ��Ǐ�?����]�z����1�Z����o��oL�w8����;�UEk�V{�&(j�VjS��U{�ֈQ�FԮ�{��#v�A�M�o�?�?~庒��:�s��q�}����c���IE��94�D��pxs�;$���/^
-=Զ*��  ?�y������odv}N^uǰ��D�Q������t����6�Aaء_队n��j��C��ֆ$j5���B�/W.�lK_��>�b�3"���U����4^�X�����6.��d}r��F;�"Q �S�#>��pa*-b�M6Ͻ�qӓ����*g�-�j�	�z�z;�-�]��f5>q�7�3����63ʛj�~"v��2'�N�#�S��Tz[U��(HP�G�x{vUr������&vC��1��}7����J�X��UTkF�M��(#���&8�Uu���x���FL�s&P���:�S���.y AOʟm�'����\f�6ੋ��&l��U�OHH�ta]1p#�{qqExf�Ϣ�x�M�S�v�~mc��tf.s�9v���O�pkEY��թU�U:����;����l[��5v����շ�O��*�]:��j�J�W����5��~������G�:���IPq�eҾ��v����
;��cqH9�N$8��"s\/�bSt���/[����.&��z��J�f�%b4����}/咸��?2Z���0gIJ2I7;�:Z`��`�n��z��s��~绹��X<�V�5K��)��i����zLez�u�	 ����<;H�G����L�k����zJp����
�?�~z�7,%���V����MxVXe���-��r�Io�r��|�8��qt |>7��'�Ɛ�jB�]�́)u�]2���S��ka�S��@RZ�a�)�B���=���2nޟ�L�C�ǭnH�B�>�g��G�H� ������0��o̩���f?��C8��<_26 �2��=q�zZ�^�-r�~I *�����O�l�K�N��E
Z�'m��~���z��Ŋ����և�zT�"Z1EOG^��X�H\5�Y�=�b:��|J)  �vq|��Sx���b8ك��V���̰3���a��d�د�����ٹ���V$��|q�-;��zRhtm�m����ۙ.�	l��k�'}�"����f�U���}��O1џ�ܳ5Dunơ��5�$�.�����bQ)Y�	`7J����P�YT�"j�߮ƿo�$ͮ �V�����H�E����H�I^�\��
��:����{u�d���xNS�	D$�6E��x�؍��r�����5�M�NN�x��{Q��@�%_�=��R.��{|���SѱElZ��/���=֖��L��g����'u��S�Ey�G�}wNj�|sK!�X"
nт<\^�����#� ��l��֙i��NKQ}lj�����a�V�G��w�� �7�$A�Ilټ���v*/��6�|K�,��Y3�;��D�smGs9`�̲�Kԅ�Ι��A�Gɩ�}CC+К����u*�4�҄�c"�i������������	�5���_��u����:7ƪ�?���@�O]T�"��|����cٽ�Qn������V��Y~���h%���5��e��T-���g�8���R���7/�6�(���48��C{��?��6��&g+z9�x���lU���1���Fq�W�;i�$֔h�;��>�\��_:�<xJE��X�9�Z�6%+�	�Afw��I+ ���'ƞ�����%�ԯ�ߡ�^:_���Թg1Kx�H�&6*v�Eސ����䣱���F�m��AY���!Y`����<�O+���+�����)��"���	��꟒�y�����f���xFN��]B^�n|TZ[�gi�\< �����ù����'E�l���e��@o`�\3}ߐ�qv��p�6C��ɓ�%�S@N�Y���(8�zvK��q�>;Z$/�d!��g<]C����A�}R��H�í�ל�,12@����~�3�l{p�vod��(�[yzl��,�i��4�1�79yxyiLQW��YkT)y�^�!����M��Y+�/�����O|Y�;�7�LrY���ø�\|�Q�V:�v��,׬�\��?wT�ٕ|E˕J2���P4`���~b������S�[�w��S+�#��P�o�O�:��IJ�����M�a��i"�l��:�mS�G2�C|��F��:��\o>�
��w����?�L_�����-qRIBPA\���|�̶x�D��pD��ͻ��CE�H�~�o�C���٢��0��~��q� EM��k��_Tz�ӂ���5��<��R`�j�8~��ECq�v6�L�r4�r�,�M���ە�����F�c�G����E��}�
��Jŉ�����
�� '��7h�]��ڿ�1D�j����ע*�t9<9L�k�[WU����i%�gf����֒Ty;9�@n��3��/�h��,�L"�Dˠ��SǤ2�p�O��K�'%P�������9���H�ӗ��Ԝ!��>�����a}�i�k�|_��Di���̓--��s���D��|�p��0����t3��)�����%�8�(��l��o�k ���Cԧ��v�A:��ߍߏ׋��L����ψ�|�.pBȂm5eN3@aYF�X��VW�3�L��c]+��N�Ow��GFFt9Rrr����-��7�l�ޓ1�^��0G=�K$7���m�_��sm$�ۣ������ttm�^.��}�2�/�s
�!S�)���iU֠G���f�֚�;�ĸE~�Ͷf;�-���xST7�+�ps��v+1�9E��g�M�+MU�MY�C����x)3:��FU�L�|�C��z��.zG5H��!,�D=ۯ�-&���wl�����;�<m���rS������ؼ�w�y�'�+<vU��S���_pd(���Y�V�&	e�ƭ�F��ubl4g�
��k�,l?:�}l$�	�+��eŅV�^��2����ǁ٧�]�C��0��1��)���$�^�={���[�s4�v���=�珌����cr̷�4yu�����,�P��Q��b����;���p�B��3��&�l�[�r�z��t�ڷ5omi��Xp��8E���������m{�Q�XF�Ɩ�/j��bkm?�_���H�z�i�f�f�C+®�p�U�蛙�����x6/4ڹvv3�^/>RKX��� D�}q-w-X��t��8��j�������9� )��+���8p�hCS��͛�>�s�FD$l���8�a�]8�(�o�5�U�u���4��_���3,��U���&�����oWw4��N�tO�ә>�C��y��-nP���)W�+ڡ|[\ ��<V����37Hl�:��Kvt�+�������?d�y��_�!�@�I�d ���ח��ںl�뛡�h�=66���h���ui7UD���E�l����2�<y�B}MN�9_ֳ��E���1sUy��u�kA�/��wSVV�� 6̙���}����QTe�g\���0&�@D��S\������ф����o�fc:	��_[3�=J뗊XB1����[��Y�nO�.�.v�_��;��N�-�#��� �H��\���}������\���%���Qt�"A��5^���=��1?Q�>}���Y"q���W��d-�\����P�9W���B�TO�Z�_:&�8�񓑣�p{�w,cQ�=��#XP�H�FL|�)S�ESG��;H��(Qf�mJ�	B."�k�U=`�b�z�N#�ڹ�&�m�:���b�4��!�_{н}�L���j�#Nu��a���}5J�����x@"4�sk�Hs����ʨ�k�l��Դ�4=��\:���0���ep"�wR݀�H`�Z��;2��p����z76]A�_f������ص�!߀"�"W��󂟋�I���U������y�ähQ�3�L�r�J� �2�����R9��n`���/v�E ������s3tn��9��چfu͂�:���[Y��/*�_���<�3�a��3����4#u�֓"��ɸ��!��*�7Z�.z�L\����]{����;��x���E'`�����\c��`=��sb�A"��������&G����V��^3�wϹ�9��.�|�kv�c_n?=��E�Ӣu>�բLǔc��z���T����qe�"c����J�E�F���-�H�j�U�oZ��*�5^��M9ݺ��bz	Ķ���w'�CY�IƳ�� w=�Zd�I�V4u��^A��� �� U�	�-�O������*����P%�(���$<<˒��d�VN�M�9=z#$��?��x'X����.�\Қ��gY-hb$%������]��f�����X3�e��"��nR����C�,��I[�>\F;�p�`��ዾ�v;��řn���w|޲x�7���������4w�����O�j<���n��I_���Uk��)�}��!��'�!����b9Z��������$�r�'9�w+Q��?�����b�`�)�M�;��Xyx�<[��{��^9�➒2�D+�s<��U#{co���U��,G_�Ikz��Bë����	��j�:BL���%
a͗>R�tUd�yʥuGT<�Y+��r>TR����"qq~Y�FB�qff�>����-�Cc�c��y^N��⻯��)��,�_����ӈ�Cο��{묡�^���J�b'7��?��s�ʼ�X��u�����.;\IU��gK�J�e��@ǫ�����%/X{�E�v4�R��&*�S5h��P�؟ۀ���ք ����;��7{�.��M<0k��+b�6)��$�k�!���o���M�}��l�):�ߐ���x���f5����{�{�n����0�1"bm���q��Bch`��uPW�WSt禔�aս��7�>�~NM�)�2{R��s}�`���j���1��^9�q�2����%2<�mɘcuG`�H���tNً�JR�]wO��i��KM�8������_�uK�j�XG�'"�J1��.|��K�������@a�g��b�V	��S$	����@c����KA���F�m���d��'lB��
�@�`-du��T��(���mb����g�@Y�B��~9�@j��� �$�.u|Q�v(u6�/-�p�P�Y��K��J�NTD
�@5�^ǿ�,�3Ȝ�1`؁��gh���]��z�����o��՘ 訃������f)
9���"E�eh�"��=I�r�N.!A����O�Ν�AW����B���H��=�͈���:C�����g�i��/����^��o��A�D�#�Bt��+7PoTxD�I�f�MTdue��+Bq�sVO����0� ���/��|�fx!�QP��!��V���z�OE��}Esˮ������F�gO�U�]��~��� �׬m2��C֠Ө������ɲ2.R� ��Jw�]y�r
����=�+_��o��	]�!��,�iƶ8����k��{S�JS�?~ة�3�}�D���JT�!E�1ALͨ���{���❳+T��Y�̘~���#��x����&'�R-U�@�ĥ��i*OvL�Ou�Rͭ���^m�R��j[T�.�؊&�!�yl�ìO�RC�l�B�y邪Z K�+A�5K|�E�>�ԩO��*��G鱴�t��P�RQ�,�XMY�#ݒ�q���Յ�����a��zr���ȈW��4!β����lM�y��8�B��Z�5S�`�^1Q�CU(V.�] �D���[jdi�O�$1zw��Nʟ9W��t�����6.cU	dt^_w��:`�|M ���!�K�ۓ�-�K���>3��3����~����*�����T���i-Q	�:9Y��#Sq	�{�8�̤
������"t:?s�m��s]�0���i�?Bc��
.��Դ�\��i��Ϥ�ܫI��=Q`���AT*S�ő�'�:��O,bOQ� @�<v�d�8R�tΨ�f�A(�mA�|�>���J�RS�N�JV/��2A�T��қ[��}��/Ĳd��aJ<��s���]Dx}vD�P��J��u�"�RN��U���g'0�#��`5�~�l/J=�l���i.�`���J���d����՜L�+��ҏ����J:��x
x�)�^M����r%��������'�c�K99������lm�ճ6�-i��ӭk혚jiJ��y����ځ�i0u2�wv�`Ϯ�f�
��������߰�{���`����Ü��T�
�ϯ�>g���a%0X����4����x�ʬ4Y��Մz������R~*�$@���o����
v-�2-�6��-!�v!g3tY�-ޗ���H'I	��T:=[����5v=}}���(SS5bT/��D`(���20j�\zx��&ہ��Ƙ!�c.U�.�1�	���2m�z����8�乿�mN̂"�ZyR�S�jK��]��?��Q�}�Y��D�>�=�1��>���N��B�)S�:�hP�D�Y]��ff�aR�p�&Qx�܌��qۯ�����tш���B]כ��6��<v�!��W�Đ��|\Rx9���{�� �� �t\�n	�K����&ʧ��,>��5=&䵲��n=h��30��,۸̰^�=�@�W��>�3�1���c��n�s�X�)��VI$����ԛ�%_�E�O
,S�ή�Jg��aW�GE"��2(���N����ݫ,���_[�O�uC����7�Д�E�ڙ~�c�i��(�Ӝ��
{��RK�+��]�Z�r=����43ui�2��|��L��"%��A#�r��{Ͷ��[��~������e\?g���fҖ6@D��~�Ŏ�n���c�.jmm]4A����Te���K���8�V9i���x�;߽�|��lb��oS��N�@le|��.�^�8�se���!<V�6����$����"��O�#5�I�`�_i����?c#a���M��u��t] iFf��y��MbdtN����������o�m<��
��|5��*�Q�~�3�Wvk�)����h�>�.2�[ �V�pq	��a>��z������a�3�os�˴����|E^���rk��ڇ� .�迚�ΟH;(a��'�#���@OR����,�vO'��~���z,�B5C� �M������E�JNk���H`~!�N��G�m���X��m񑕤�%��gp_�����-�JBT���$��ieX6�c��(\L�r݋����bn��]�#i���K�ʷm���eRq�h]�^AF���a�����FK����=�-�j�׎���ʠn|���>bH(�����"):��qz�LA��)
���%w�4?�n�:⥇��*�XYK�4�j���ߝ�
�^d��Xq-�߫J�p<��I�u˩�r{Z.��9"zO��Y��(1-X��Ø8��:{���Vs����P\�M����Q@No{r��g¦�ڄ��t���VZ)��v$/�f��-}�,����}�a=��e�f:qռT�1y�+j�
����s��Q����򕋖�����}'��36�"���b�ġ��gjieGF�A�D����wI��ʓ脶�7��F2!6�����1�=2p������MpetR�����Hcߝx����K��88.� 3�wY�����b�����r��(A|��j"_H�ڔT�#ΪNˤ���rhB���B�lB�	J)KE�h>h'�f畱�:0�}��Ve�2Jy�������r�,�.'(nS�. G����01HP$����Ι��:�Gb������ހ ���N��3�¸\y��|���0�d'β�;�5Zv����b݊�/-e\��[{�/����UxZlyUT���g����V��d�we��1,�1t@��fO�N�fV����`e�Y��Zs�A����彰1F�a�Ɗ���?���m�?:��B[$1�d��Y���_��ʾ�kfvy$��c>����������R�O�$j�o�4oj}T>.9<�����PUk\�\��͛��U:���.�O���"�6�5�i��a���u��.�����)��t�2���XI�[���=;�JI_�'_ck�i��)M� ݓ�),��x��W��B�*�S�k�MJ�n�����~*rg���rT(8�JڣOݟ9a�s56�v{dWR�ɪ(��A�g����`�A��P�=�=�����B�-e��1N�}�o�z�!���y�՗T�%���1t9?��"�-��Eg��w��R7k�.��O�Cͽ[�gȗ��/.�f�O�h�y��h͕j)\;@ø���U�3���Y���N���7�;zb��{�"�YSEDṋo!QѪE��ª�v���Y�	U����}���?9���BP�����g\C���h\�_l�mi^����ǯ��|T`��"R�7H�n��~�C[��V�O����S�9;��\�ay�Ji�P�A�A�+M���z��,�ClC����2֮���㑢���|o�v��!G3�岃ܸ���a=w�����@�2+;����L8ݢ�I5�ݸ)1�@�F��u�R��:�U�����O���ѹJ~Q��l���ſ��vw�ª��̮�Vi&�L���M�>x$�s�A�U��#vE�܌;�~�d�y�k�s���}�z�����;LJ[o�����p���ߍI�PT��Д�Hܤ� 4gg����Yh�e�rF�"�����`��D4*Yh�q��t�N*�|\��y��bΘ�R[��6衠�5��&�P�2����4��f��1=G�/Q�m(�@�wR�I2��$:�~^+C�_�,@�nc�3�����7��xq
��I �i�|
�o,c�I�%�s{���ʲ��ky1����S�Tj�Ӗ@Oj0u�Y���4�{B��Hw��/�l2�qߙe !Gg��K���u�Y%�Y���ȗ!��؊�M �/�	S�T�`n�U*�栰�T�@�>iſ	=��S_as��!r� Pvaw��fr��N�z�<��P%���~��#��<�n
=ZD��&z������cC.s�T́ϑi4��I�%�Ȕ�5��5�p*_;��^�A����D�*TJ�:Sl
TJ���x2�!㇀��c��>C����V����
�.�=d�}��a	��q�xI�y����<���}�U>�rn��k;�����~�;����t�C~��Q�833�`r��b�F�W�Mr,e�ܗ��W^}�;� M�ܗe
�eĿ7��uP�bI��� C��>̻��Ox�w.f?�@������Wb2P^�d0��3��A���m=�S��j��c�.V���8�� T���#�lA��l����G�s����Z��a�]�9�m��ѡ����$��P�٩&cb��F�-��}��%i�|g�*Rj�!���ͱL�~;�����jh�Tx�-n�q'.�n��V'�P�Q��In�R����biC����A��}bF��.?PG��q���K)T��Mg>�����ǩu�QIn�3��Y�~!�q��`��S��:X3�,3uqt9fs�Y�B��"6q�������*_E�N�קg���m?�i�5�d�X�oX&b�f����3SD�����Ҕq5!�8!o��ˢ*�)��*.Y�-2%{�fd"w ��pf�(}��o��Ê0װ�w�-�S�h�e�^I�=%���`R@��|%�~vP�u�;�&�1Nhg����_�uPѾ嫞%���ع>[(��@�ʠ�->R޸�R�Ǥ���"Җ[����dW���3�5F�.�͗",����v#�t(*kR�]�b9�O�洔�"��O$�Hh��[o�v��f�K���M���5͙D$cl����p��:��J/5���h����eV�K�������YRrN}M�{��~&���TKc�V:���mIh���^��V�VDn�64�e��(���X幕���Fzz��o��OP�E9lֳ)l�4�h����d?]ꟶ�<&�H�%x2��Qq�B_���	D+9l�,�^����ߌ�*ήk��'�#x�{y����PMV�����We���_�W��H�Gr @��I�}ʏ���D�|�4�J�v��#Ȧ3'�xpv�#���4d�������$B���L�\k��u�Y0~=� �*�і��1t���Z��JV}�q�M.���EF����s�p�:|��c�:�H[C���ڡ��J��+����v���k�w8�8����(�7D�f��V�t�����j�)��l����׺�^�U�?�Ȇ�҂���%lg�.�آ����j�9�����q��2U6���m���I�V U�Lp)ͺ��o͙;�
Y��:�m+����}-0�ճ7r�h�'������aH�ѱ1�Iy��{���]�]U�0zs��͔o'���qz��v��S*�3�YO߰mϊ�z���%��5�9����9���F���Ϛr�s�����B\0�V�ޘD����R�H�l��=p3k4%��,L �ba\�qp����}^ݟ���۞�eA�[Jc?��m���Kա6�~��*�S�^\� ���K�~�S����W�'fe���l��Dtk��J��K��\c� C|��x�QX�cW�F#���?�^Plo�s��*�٢�77 H��I��*nh0׈��E�-��w�F�m.��P�wax��9E��ĺrD4���$�gZ 9t������ʀ��l�c<K�4&�<@`�M���d�,�hS?y�=2��wƃM_{�&�j3�!��5��'U=W}j�
�I�T��,���}�n~�8�����ʓyW����7��΃Vm��p+���L��:oΔL�1�m���`"�m���]����~�)b�ȹд�����:y���ɩī� '����]�y�"sѲa��+��u�]�^���C���&9����<��<���x6��ٯ��'�&�DmĜ�"4�9�%�S��o��,`��pz��/�3�K���}ᘘ��V'�l�Ф� �cf�:��B�$E`�>�gP�Bz5R �s����i�b�����v�S�@���H��A.��4Q�4Ez��D�N��包N�*I/"����k!��޴T(�Fí����14�F�0�(�	I2�q�~���^��^���h��VP��ьW�ᦕQ�E�Tӣ
Y筯KK�.�$D�W�gp��Q~ߺ���z����<��8�sV�V�Z���t`Va�U�F�B~7f+�����bi��byD2�9���I���Q�5/L�r�P�dyՌ�h����Qk���}.�u�	�[����%PD�BQ���LV.�����)|��U�5/!������\ +�+��������2A]����]�>VeR�r�.5k����A4��daw������kN�fI��ې�)ꬑ_Z�C����]ύ��`UN��uqڥ���'/���\�8�&U_�ȷ�A<K�����ǟ�%o(D=v�\��l]^u^z}��A]5Aa�T`��0���.��w,H�8w:�<~hM�:v��O�k��*T��1�klQ�J���n�h��{���ˆ!���,��ި�Q���i�j���f�\�]����Hg�Ce+0�_K��Y�m`�f!˔n~�'OO�*O{2��3�|k�Б��(>(+���c�������C!�j�^C�a��_@$�f��޿>^���)s��i����ÛH^���}M�2�-kg�����Ŧ��oB=:)O��񕇚5�L�hwH*����V�{��n��h��ٳ~�#C�ȗ4��u]ǰ�b��q�-�Z���UyaI`Aq��c���>�5�c({�IqehV��[o��9`�fl��˪P͠6�����̛�g�E�{*�N̄���D(U�\#I@z��� ���J�y��-]�-���#�� Jy���j�mYs3 �?�d�$b��F
�Y�K��R��S�%%�Q��t���rL6FKt�DCՋ�("��Y�#�i��?�����ޥ���sY�L� �('%�a?�q����,~��AN>�w�=s�A���~�����.��K��dc�z�b�͖����A?:�z���ё�߂	\���ξHF���^L�����]hXb0V`Y�bn�[�Қ��7q�r"h�" ���_�d��`L;}���qT[w��8ԇ2�����_�w��,>��&j[���J�"��x��� �p�Y�T�c��75�~�~1���X|�_������hd�f��-v�K^�8x�L|��ϒ�b`V�z��)

���d�<��"�E��.J�r�H=���/!����j��NN���-*ڝ)�G����Nq��:���������x 3��&Z��RL�;�4�F���l�0��U�>��l�kFy.�������t�p���Z��=�?�*��D
��:�M�rt�=�~i��&0ԏ�
����0S�o����Z������T�!�3�`Ei ~�H
���^O¯�8jg�����s��\ܯ�:�5E�T"r�:_����w<ś@������\<<;���냓Lr����~#NΑT�,��T�mO֫�;�_9p�\�.X���+8�;�UMf���m���^��*TY�V_Ζ$Ҋ���}�z��!��~�KÕ![��6���;w9'�����\�� b��o^!��ߵ?��5.�6��/��s�>	�Sd�����9��j�����W�����	�
�c�G
�=R�>��.��@X`��|����(Y[o��58���̑���#��@� ��?�,0�Hہx���7;�.0�j���ɬ}Z�"��77Cx��I_�V��RU�Jj�������̌�-W���\�F"��O��yG�a�����V��ց����#���r��5SBڧ[����1T�E!�FjtH�����j�ݿ�ۡ�A��t�v������wώs���.��/\�f�I"��bfg?d����嘵� @������G*�"���P�>�Z�
82��zS	FF����L�'eS�5z��4c߻3�5�}؍�s�u��cg��2+�G�q3f�+�����o[�M�8�f���4���p�$8ໃ��nn�\�h�|�`�dc(��B3�����1���`�k��������y������Ƒ��3�\�zq�5��c�s�rr:.V?R"z%ރ>��`�s���%D��֧܎�LGK�*堃������0d"f�'I#*�$�����8Ɏ���p|3����P�X8�1����Z��jf�ǥ�(���+��ֽ�hҖ���VzIN��[��b�Ԥ1-�I�?Z��v�?jm� �����������,������K���P������(�9�Az�@�t�U
U(��kc�
�D=�gS^L1��
�f�,	��գFm͋	e�q+�h۪V��z�X���(���^�����m�����)��^�Ө"s�bn���ɲ>�w.�MX�ס��8�
!��x]��>�
�$�;qGOj�+�?F@@��s��*����3���{��)��7�g?�G]z	=j��3C:8�~��ހ��jG ��/M\�m+a{`�~�a��]��&(0>�w}-�n+��OY�	�6�����K�r�!Ny�E��9��I3$(��}�<�x�eD�7�����X�g�Xz��)�8-�L$]��g��8�C���%>����I1t��Y����0����h�Դ�����qp��`zfU��qԅ���M�l��q�_�bi�tTp:p�{��xz�Z|�nrK޽qh�c�q5���<}��p�f-��|��ڜK�xھ�D`x~����\�DWy:Kpd��⏜]ԗp�T|�����(�=3��S���{���_}�}id�)��)m`����1����y�c���~IA� �����z��u<�����=a#gqe��Nk��59�35�4L��uoɅ�F���o:����aRCw��V��뗩O��:�p6s���;��N�%C�U�KH����SJ�J�K�M��KH�io�T�^!�7�$������ZSW@3�5
K� E���.����,),at�\��m�\��������{d�}wƀ��]/-������P0ۮe��i�D��׿O�֑��W�r9<�7ѭ��
8��0�����"ɍe���'�x��Q%�9���i�N����@wX�rR�O��1�E�� ���^�1�����rN.x�����TM����P�_=&����W��k���wl&|��F	����ڻ����m:}h}P���V����=� �Y��Xd�o;-F����	�G1�4mh�;��b�8�����cjK��A��|n�YCi��KH�ї��P��%�W ;˯p�lDp͕)��2:$uH�-y�}�Ѿ��͙ٽ�ɗ��[װ�o�Ţ��l�M�n�����[J��o������x���F���7!_�s��7?���]��E�Y�`�}
y�*&��[�E"��{�^�k?o�RUsn���Ph�6����90��q��(݃4���A��_�b��{�z�3��C��opג���ís)ԙ-=�2��`�����[�T��;��"��S����MM.����夰����^�
�`ߚ4�}�y��W����L�Ge�U����x�z���Z6�ozCH�br�����m�	�ӌZ�qM�eI3�	y��:E�oWH�;������L�7[����HނcMSS,�^��:s�N��l3�ݑ@�7��a����!���Vu�4N�A��]U���IӨ�M�Fs�����("����i�m���P@c��b�}4�c|����Faiˇ���@��U:�1T\Ԫy|�=)���\�eK�z��ݤ"���%�������99��0<�e�%�y�S�,�)A9�0�P��8��Z��b�{�Mg�����J�_¯y�f��m��c��+�	��h�.��@-/omS�(�3�F�C���CY��j��y;����{b=р+A��CEQw���8�g-\��UN��y�OT8|oW4S'm�79͔�����{�I���jkk4����
��ǧ��2�Cm�[�
�B�����d�o�|��Yk8��\_��s�sq�Cgl`�h�TSU�u&b9�d��7İP���9T���&�z��7�  w(��[ړņ�=ؠ�� ����F���=yG��$]m�w*4��~N��z�m(��ӷ�ttDö��%����ۛ�Yі���|�ʹ�ɖK����H�3I��PZ'c�|�Q&��6���\H)'�=��Wr��Y�ߓiŮ��[�r����=��B
�gXC:�mEl���3˝9{�/�����]k�dD2���k��˓�Z��O��h���ƿZ������	8Y�Z塻Zž������O4Io}}�	���6	l��h���#����S.H�?���k�/k�>�k��bއ|���.�h6���L+�#���s�cZ�׷�qK&��ә+��R�Zzz�'���~���^V�I��W�+p��Nu�n��.^����;��g#��vVP�x��}�F� �. g��ƪ�F�D9լ���65��v���]�_c��&���a��[p!��[`<�I�
B���gh� =���}�G3�ǲr���]��t��թ9kL�y�ou�_�����[�fu��ͥ@4�Z���+��{6�4�{x�b5�o����Fi�{:����7?��B��{���Tp2?�0y��蛈�2�"�� ���رB�6�ܲ��.5������6>�i1���*�0���WH�F��Y���p&���v��TfJ7hTb�y'��g�,�PX�	䀫[�c�lvl�F^����>i�x��8\�R�����kq��Z?��d��eX���u �d���u��;�V�y��[��`�"h��i]����M�d��/�z��/��@�_��e\�	��~��JWO���:���㓖�3�:&�J�S)�bL�� /Ϊ��~��R�����r�ͥYGL�����eF�`²��[����'��<�|YYY��g<K<����«3�D��0����5���σb(�yĝ ˘�ZE�����V����!l��+~�����Z����SZ�N_��}P�Ԙ�[��k+RŒ`V%���p��)*�=�|��$5��!5\��}��2�nz��J3�g�>��L�q���?sI^_�c��F=kȀԹ�x6���֜E�@	���8��@G����1����~�I�H'��j/�_�Uig41���A�����5K$�Na��?~P������r�)���z���^�[���^�	'u�G2�y�v,H���T��p�E�3'���1�����*e�TR�cOl��'�{\ٯb)�~�[�O lk܁'���m9e���2��7�Qڌ�"U(�+�%"��ص�`PT\|��W��B�F
`��詠]c��pi�';�o�|����z�qHo%v��@0�r$�����>�J���f�/�3;�&֘f�=B�B�k��)�Ϯа��C�u�5��<�Jj��.�#}�4JO��h�+���D�c��<��B����z��Z���1'"��F�a�+�~��&��V=�֧��AX=P���Ͽ٩���v����L����z˨6ڨ]'�KqZ(nmqwH-P,��ww��-(�)P�KpR������u��+kM����ޗ���{й��)ƅ*�H�'
��ڥā���m��Ϸ�� ,��^�<�^�M��8	��U�0���}�O[���a�el\h;���\.Ӵd�@���%Q_���?�Y��Ђ�	������Y��~>>4>_��6�t�S�����`O���?��X2�㰹0���c��
ި�m��ױɱ�x,�r�{]+�-(���)���\Q�r�n��
�xB뱙����r�fΫ�0_ި�ϓK9!�
Ǥ�m�H����=���62�~t-�엎�i׾O��্���6��5cݗ�G���[�hFV�	\kRca��&��\zg���Y��Fm��ZgM�������aO��ѿ{�/Ckz~�/�_�ϼWF:@�:|�K�E�$[�ꫀ��bҤ��O�����v}iEY���:g�PJ`<�qu�L�#d�Ӂ6n�M1㩔�ٯ���K����_��N��dDc�&�C�C��i�ؕ���Ù&�_�Oܒ�/��,�s;z��1�Յ����ӻ+�V��k�{�fv>�wzGn{~s5�4�G�Y6.փ8�弩�%[А���Ry}0_��ڶ6|40:��1��V�̪��Z�e��j�m��b�fj���W�2�����X�����P�?�]������ZH*&PP:^����#O���T�B�w���6���j���}�CJJ���e����	<Td��2i�P��1�Tq�Z ik�j�R2"���	4$�۶�6}����U�.�D�+.ޣ�k��~� m���#�֌��7�íD�Zo���	;�1H��Q?^ �g��r8��o��]�C�K��(gnߥHq���^9��]�$��戥�I*��E�:$�/�'A��@� wD��#�g�z�}
����K-]���W+Nӗ�+��2��6[���;�YY�?H���>���>a�(3�G��D�efe�
�mHQ��)���3x��1nE'.�����Syx��f�I�@�\�2�b�����W|��a�;�Xs��_� ��,/��`_�8Y�y���@����� u��������ď~!I�9Vv��^<���O�����'ڇ<�RQB���^�i�q*B��d���A��[ѮK�Wk�B9�A��G�S��?���x�
���}�o���.�����D�CRE�F��WI�"c�����8���jZ_���������,s�9'v3u��Xk�E�7���S��71��J��4��[\��n���[��ЬOx*È����+mǇ�JTC�朣|�;{ǝ�x ���%�,�8q;X\z`�x�,Y��
J�N��$��X�#�I����VJ���(�B�V�Y�&@�{n�hΖ��I�K�����Y�׾�
�Ġ�bո����ۑw����}<r6)	_��?!��&�=�9�\�,6p�`�m�����VR�TM����`<��K��p�尾�}�,~k�t�<�����na�q���P�b�EI��}&l���Y�+?�x�]�97�;G!��q&߬��	K���_*�߰����k�V�7�W�88�F��'��yc@LѥJ���E��++	v���17y¦�%�h�������y��:�����t��M�B�YS1��Iů�t��x������ 2�,�槬:�c-��@�yӲ�t����[�����ǭ!�n�p"P���fh�^,w{��ah���;�V��&_��*��^����G�49S�v�,f�~� ���S���h.�\m��Z*����Ù`�\F�)�U�*�*�[�`m�%���+l�����al���� �e�{s��'�fK�MLbr��_�U2 Clc�,RBiiis�j�PɎ
���eA�0��'��i��r�9ub~qb�7��>��=,��a�j�wH0|��kt��KKTV�hE��T����i�M�3:���ɭ��ᰛX�ji�=�v0�a�%N0.8)�}�1��Y�\$�5�wL�dvb��٬�$�C۔ɉ2~��v���M��Cw�!��v?���i�j��vf��V����\�v&ILX�&�$C�~^�52�@?�����E��Ա�-�!Grz�9M3Ͳaq��X��O��If"��Gΰ���O��<f徧˂�>\�����}8{���Z?��Ix4W���_V��'�n��k���"|Y:��wŪ_1����A�3�a��6�e
��O�8�W#	W�<2�����g�}��`���E���D���E���5�:�&�F^�j�L�����H�^���r�}��;����P��1J�^���Ccll4d�0v��Y9���ڷ�왿��6�0,F���Qɸ��;U6"B�w�"PY#M*H��Y�3F�"���@�]Jn�?	$��E��LZ9tK��:��ڃ94�Ƽi�܈C1��s˭]�Q�4Ș~������i���9�������E7Y��v�i�6�L�2����SG���(���-��:�j���*�a�M�ߙ��d�P��ׯ��),vKT���z�	p;Z�����K��(�9�*eM�_c&��1ǢG��S��m��<�r�3p`P1=�k�\�{t��bȝ�JK��[��sVߟ��s�u���NNTη�����Fs�w����8I�L�e��_l3� p��&0^�*-)5S��4A{�S97�'a�9���&�#���ǳKh���4���C��i�۶��։�@%Z�������6`L}�bZ����c�m���ծ\6�L�#/�Lja�/?��\�|�R��N�=m�*2`f��m�}���llm����l��`�r���K��Q�]��v��{�Nۨ���q�׊��q���������S_��C7�	��ٺ_���:\�Tvghs�8�+��F��#^����;_����鷩��XH־Cݮ�u���C�}�m|n��]��=4������ˇڳ�� �Tb)��u�8�G�YzE"�G�Y]����:�g_<�����7a�V=�yo81�U(�-��ˇHn�L��;���	df��W�"��2�4DQ$\�V�L!4���NSj���B��s�OS���L_�A��\m�;o�; w�٠<K�x�?�NMg�e�tdt����W�s���Z�f�\R� �`�����&�<I��-��}����w �2�:���7.h��3l���<�����>q�_`���v]�0��W�6Jpc"&8�\�*K�%5iߥ#�*�[1�N�瑱
�^����w��T��՜c�^n�����L-!�禕����n�ēi����<�.u7L`d�&�J����������P�6�g�U�Ƹ凓�q��Vjx<��T��v1�޲t�_�KI 7�$�J[��D���&��9�(NQ`�]�/I���s'�������,�E)i��;�T��C���(���b�F��O@�^�F�c���������`��c����y�sx^�<�r��_᧩���E�{"���D�:ѫ0�Ŗo��k�G����� Ѯ'�Փ�lUޟ�i��:7o���;�;�����KY���BCo:�����&�_�I��Ì�lF6.#m�/˧W~Sϲ�I���J6����@נm���g�C��[%Վm�pv%��6�� �\Wd�Ϲ�'�p�NX|�$]O�J��1�����Y�w� ���s���R�S=��I�/��@�ɞyz����[�܂�.��B��D�1Y�Ȥ럩���}*�ڜ�|��<�~��A���7��֌��y<+5XԿn[k�b��P����ﮋC?�~�n���i�&�Z����_���$4�Hq�>|��P���TJ��Z-x����e���gQ�4S�L:�@�H��C2�@��У*���w]"�K!@�YZ2dF#�|�ֿA��,%�㕑Q�VG�t�V�~b�ߙ1z�w�'k1)������e��f�j�]�4��}c�����t����o�o����|N�iWG��j���}.���W^����(e����;�L�o 	-��1kC.o���>�:�\cef���_3���D��������Ox�:]��M�����ņ~niv�[_Tݜ%;��9J��;���Im!u����sQ����:���.ܕ¹�kTj�n罊�;���Gv�[���=Y)g('��zCy���p9YE��1���lmo7���edf�r�j[ �Ο��wt�c��6;= l��M��81�O(eQ!^���z��x�` gr(����{γ/���&56g�0�������]-��y'�ս�������E��:��7�{�P�Q�L�b�,;�p�	7��_^���"�*�ޟ���y�$���W��ߺ�ˮ�\y�۷��7ޤdd��Kr�o1��i7�U�� .E�?/y\G"�_G����������wz[~�I/\ Ύdֹ�k}��]?�kq�����XGp�������\Ư������dI5��N�S4�� �'�NPUu�����wx�rp\�̞��Q�=�/��?��<�"[��\��RT�cC��rn��^�<���AU ��'f/J1eK�W�4W�`3��|��S&X��<�<��?{~����YCyo�2��)�U*���D�\�kh��lp�S'�x��ʮ�i��yД:��[8���׃8lP�n*-N�틠֧���4^��ጅ�jJ�t��İ�+8�|�$>���م��JW���U�W6uӬ�
��ݴ�r��l��R2�E��IfF?q�o_�r�F�t��?!y��l�$���J��i�M�o*��e�R�l����M`5]�6���ٖ�-G��B�0�M`c�]�4Z��xKz/�BRI�AE)U��%;���h���QW�r(�����u��giY�$&.���C���Xфe�ū����Z�l,Φ ��]%��h����ώ��� QO����U|��K�r�N?f�eS�%55т^7����ҙo�&�����WVŞ�&ns�q�=�y������>��f��lCC�b�an�J��|;����z� �(�~�4b���������ܴ����Nv>R��|i�"F������p�2=��=����fB�f吽q�۶m��sї�3F����2+��g(�ڬ��ڷ����,Ǔ��ni�����n���i�����RMM�p�zj�ᇦ���f��ۼ{u��I/ޔ�6�}m�,1�z��O�ә\s�d�2��oFk�]�
�)�zਜZ�
ǬM��+A��p�l��ala��:%�?�#?��0)O�b7���7_-�$����}�]���'PtvM�]�d�}���N�)�K�ᙽOP��Oc�^4J`�G�<�N�f�N3P�'C$�U���/CǼcX3y\Uю���Ip	�,�o��e��,�Қ�(�􈭰�|��O�4	d�_T]�1�u�%�w���FWI<+�*�ܸ���,N����H>$��+�/�f�p"p���nM�V��6�%1i�n���_�3���>�����$o���2u��u�)�[1~����l�5��l�=3���G�U��M����#��&�[���*j^(�ZO؂_c�a�P�=��,���:v�~��gi��3o���A�U�.�[_h�������ib,,��� pQ�e��-zl�K+��|g���v� �}Ş��eu���{��we��N5 �N����m�N�<���by)s��jט�Gh�rِK��8������us��i�����8�h�};+u��� �,�*�Z�).�բGѥ������Hc��g+k0��ぐ�V�ݏ�''1ݗ�Й�s���NO�,4G�����t����Z	����Qm���������Ds�p D�j�\��dU�޻�� j.���]h�)O�����9�&�5��Lχg����D�ri{��.B98Pl��A�L��S��aB�7�g�D�;=1_窈�w	V����)ZX5=�6S�\sm.N�����Z�������3F���k��bxt?qJ���g?]�Ε7�l؅ݏ�Š��p�t~�<��VQ����ླྀ����
.�6��{�nao�����;h����<!W��PT^��I� �
����q���(�Ҵ�A�F�̊��_ɷ��p�V���z<̯3|�ixllb�%��w�͖c����R�iii����x\X^��K��ap�t[$|��5f[��.���}�ac�bg����,��_��c��w�3��-�M����8z�������wȥ���[�1��������=��r�m��s��}0s}ÌY�}�W;��0��x����(
�͂pLt���Sv'���mp��.�Υ��"5h7X���G��X��vK܉y?aWͺZ5�'@��L��1���s;������ץe�M��� ���G��/�r���~�t A������F�	�V�N���mxddwѡS�cM���N�V�b\�ѼN�u�w��Ɍ����e���#G~�{�����z!���yS� wkͶ'���YhJU�f\��ꁣ��DܢW6}F���� Z
�/��0��"J��0HD�#�ה�٩�.b��a"��W���zN����N'����}��P�Y���R8�r� �9;�}I1�4����B9�iT�b��<N���h�n2�d���z_�h���D���a�e�z���b+/�IE�)+HFV	x���R�}�l�Q���E�X�V�c��Z���׿F��}f��3�?:C'��aZ��V�L�rE=rN7��u Akt� Ir���c�?�!?��H���)557n�Cȗ���?�5/�����Z�Y�BˮH"&A�;bw�/8.��B�����Tۮ�p��n�go�H�l����2��"�R�6�l3���#d��QD>�T��-���y/�}��u��-�T�4��c�䔘�k�e^���a�f�[���,ݲ!s���Km������9->��O]��пlӁj�Y��k����\[_/��`������Օg�>e��k�P�Y~f&%��ۖ��Y���d%3}�ܿ�`���>��J#:�Ly�m�m�i���������sE�����y�$�� >nNc������T{�2�4+����-d~��F��K����/ڋJ���W/?��=�Q�RWd$JKǁܐ[����;���O	�@Ic�|�������9X���@��/����K�܎F��}�6��@���M�b�T�5�H��|��<�`zZ1�돑��ߗ�����=�Pk'�T�T�$͢�!.O�!P)�>��=?_�0���o�K�#�U?��t-}}�A���ms��~�۽��va�����'���Q���s���]�F�8a�dp���W��f�Z�5�s�	��䯀����$�߰�c����%B{��6��,�wm�����<v=ϝݚ;����$씍\OA/WrF�?]��>U����&��`�O���'��h:Q����qi��ޮL��߁��a���U{˱�j���n�PĔ�z�!�aU@� ���^I��MI���󢎞l>�~[�����tm-�}�C�=�P���k$
U���n\~Vl�).g��?քt�TVV~-�6���n��ݟV�;�5�S��B��Uv�6�A9$��T���%*�}����F��w�&��Nȯ�[7��v��w�/u�;�x���]�������׉�>���֘�I��}]Z��e#OO�)h@@�/Zx��Chb��c�2�E#��	��GQ�02���	���[7������z��;���K�<n��[(o4�5=w�� �=/��\���>�!��5v\ڜ�h��j�x5y�C%%B!�_�"?r�N�>L��v�����N���HD>2�TI#�L,d��m�P��/�"��8�n�u�T�;���K�kERs �WYX�/j��|�&�q��x�yr�+u����cy�(���@]w�]���;�����-؄�������R�7�z_I�EQ>��}a�D�+���RTܿ�-ѕ�!���)���*�B�98�6��j�&���9��P-�k**l�z2�F��l��]!\����H$RxV�:�]�㙣&��U�o�1&?�I������̹������UXX�Q|N���@�q��ŉ�����@��!��t v��Թ������$��;�F�L;�qk�����Z�%D�o-���[;v�-�ג)�y���Y*��^�;��Ǟ�b3Vpgo���:��)���S9�4�A�	��*�;�n���U�'�{U�.����߲'/�5���X	l��́�w]��p�^�W��VгH�*��6]<n����;�O�;ϫdr��E3>����?�}�@3�,���bGJ ُ���+ߙHnl�\ϭ�i��k����SS�K.3f���v�k���_u��##v!F���
*�y$�t��v鴍:'+FbY&(�~�����v�!O�Ȫ�����ߞ_���sui���RzleX�L���̐�x��x��9�l���\��$l��JT,^��=���M��������z�Gnױ;���ʹ�
�A�Cj+AB#������6�˻-�M����ǅh��a��P6Mn*\���	�ƚ��8�2e#gg�C�@�s��A�Q�������y� f�U*�~���|9-��y��]�_�F$a��WŸ;�&14!�;AHJ鄂���1fa���,�_]%��<'4�~��'D�t����"j�r(������K��L$H��<�f\J+V��߲�����d��̘m��s�Ey�!��bh��(���h�������R�]?����~Jk��'!p��;��Ns#>;;�Gl_E�4���]�����ے�Jʸku�ܜ����������c��=qq�Ϲ��T����<Lf��~($ED�O3�Jg2��>0�0ю+ /���p�#J����?�Mh�bo�Xj=A�DuCF����ΰ�Ȼ?�:8�DA��گzU�.R 
�i��3�0߫����\����'<��$k�4��zKH�NO�q̃�v���Z������o����zp	��ۡ2������X��g�8������}�6 +���<�Ϛg��;�7����Ikzl�l!W�2��Jy�k�Kk�w	f�R4��W�~/������t�/ǳϴ`���JB�}>&j�+��|L��zO�}��L8'�2N�qTzڵ�*s����0�W_�o`�	�.�ޚ�\w��^\�:&�*�p�!�艠�yiԛܮfe�eXo�j��}��n>��]�;�ئv�w�
��B&w\Z#������`��H�HvK{`hW�`jO3�`�P$d�?��8[����;��RC������o��_] ��?}G5��<��P:0ۇ8D1QCQ$�PSeN�^�|�B��*W����8^���>Y��
��⨬�t|Z��&RϥÊyk���E������'��L��/q}��h__��i�s���Cm��sY�� <�t�ʹ~�e��P4p�M M��q�<�L�Ar���>���dϛc�����+���!���ݩ2*\�o�d�m{���>|��a
 ��I��r�&�K��SU|t山@ ���>kT׵�ϙ��יa���z_iWVU���.�����ĩ�t����X��B$������y�8o�vn��{m���(����z;���\^����y!󜬘�#��ਫ�w)*$0M��F��}O�����;�{w�7����w9�ک�M��WBx ZYW3ڍ�X}�ʒH&�v>n��ei5"F�@ ��fL>�U����ht���������Z�ڒČ=۹�����}�G���s��n{0n^������55�O���b6��)Hj�(�J�n���
�r��w��e�OcK�:������[7Ou~K�Y�/�B
�,�RD��-QP(t,�S?0W!
4��#�sjJ����S9���J`0�>��8BǤ�^��x {���B�I��[&�	sqt�EJ�-�o�4���������C�TBE���\�c?��q��PF�Sq�>���e1(��Q�8�DJ�"t�6����U�fF��g\�c8�x�H�n�pcO��A��7��EGs�O���D�kk3=�ۥ+��~ҏ�Z�C���m5�x7�ʰErgY|W.��Rě�	SL�@{6YP��/�ǉxߛ7���W����T��ݶ|҄} �Ϸ(�ޫ��GF�bLt[�p��[B]�vV۫K�Y��*��&����Ms���JHj_��u�^�#�]�U�6.���4�:_�����|.&��zz��9��=|�{=�����!�����v���Eq�U�����`t:G_�V�Erl���������7��x�7�l�)�4Y6�
I|��V�U���ـ�^H��= ���(�=�f},,�#��k�}��P��.x*:m-i���@�gA8�O�<w�bʹB�c>w��c�n���O��.��Z��*����F
b�2K�E�i�H��谥�zb�%�6�0G��D�b�dccͺS���ۛ���Th�7�,m$ь1�Y@D���C��=�J� ��#���<��Q �'���^ѹ׽���7����t��8-��ؒ�R��ii_о�`���)9�2��f/=������[���+���ykYM+�4@O�[��xT�5{mZ�gd�BS��7��Q�=u��@ ���4 �M5v�"��]K���UX!��[��XY� e�S���;a�H0[�U��t1��v҃G�KV�<A�~ч?o��P�9�{�?���g��-6hX�c�h'9B��P��)�%�<d��F��ZX���&�1#O�fB�%S�����߹EǱwǶh�7�]_��y	� Ox��D�r?�0��r��x��N����:.�c���p�� ��(p��b����m�zm����.JR��]�T�z������n�iSU�z��'�
����Y�Ɉ�o�DA�m�?�r)�}���ĎZ*�>N�<����7=vtx����9~�3��X4�x�$��OFq�213��ZT��#sU�V%�*�.GM2G��F�scxrFǁC�K�n�sY���-�����\�B�1��v�����1x�I�������s*��x�����lg�K#�bj���[I�E�w�^U曡m�Z*����D���Oe�Ə�}�s���v�,?$!���U���� U!�m;}eH� �(fd�-Q���>����{��Z��w!(b�,"�4TiL�G��T0��6�*�\G؂GKWT$ �B���g�O��
t(���&H��+g�9�����R9&��
�u��JBS%����1��{�Q�?	˽����שq�cP�����:�X�G~. $��"$���FZ���zk��plk �uP-~1.���x���:�����L��^�po{/�������#f�q���������6RQ�l�T�m�_��C��:*#����2��ė.<��|�����e˦񑪘�*���i�
I��
I�$��J<����C�GJ�qÿzP.:��᤭���������z�M�%%�&��MO����G'*���t�]����Kb1��Z��4�/�e.���0|b���5��V��c��D�hyg ���y��\Oѝ�:�����4�q<��ͬ�x�T9�H��jٿ�������OS!��؝jr\CrssC@P!��k]�Ȣ=A/�J�,'�9\����ݯ�y\�����b���������ر��\<�0n+�:-��2�-�Q1w,	U��D�3�ݼ���M4��T#.�����&�]�d;��K-{����OoՆ�ߓS�}1�����)"DR��E�T6��x�"�5駷�N�+9w��ȡ�E8�0#��&�f���E�HI�Y.ߝ��)���x�飐�yF�@iV�ntV�X�"�C	2���ot��d?ţ�e������7d (	A��a� Z�9��Yy>H���v��?�YE�n� D���R.a�_5���lngw�/�~�d�ĐAar����U�G5 'ߓ��] [�51�
�4%$ eXN��k륳*��/K!�]�d���ۥ @8� f�!��%�"�R�B�{�3P���3��{(I;�f�/_KG[�JQx�]ee�keャC�C7�Q��*!��X?\r����ԆK�6��,�_jIk�;���;����>���i�����)c�� H(��:CM��m�T����.��		�S��6��g�L�4�+���H���#?���<��l��7��7�_�/}�t�w��ƾ�.���|JUr��4Z�ΉPS��p�|��� Y-ý)��@N����wc(��>�O����|������C�0�~b�D��hyР�PRc�/�L�v6Н����gw��%@=s���S��:��� �6R14���2��nWzj���)y��T���]�l�A��Px&g�5*Z�`.cC�7�Ū��$|3:;8H�_���Iz��+�a��2{e>��V�e���p���W�$X�MY�����������z�Ҿ�-�S�%�{�N���b��o��q���o�z�@	��M��?]�_�r�u<vl`Qe��1�=dkB>�Fi�;`{:�����e�k~��@�S,�M8u�m�ð,�������b�`��=�C7�hc��*�]g�|'��{��K8~���*�>rŠ���ؗ?X�[�R�)�%��7�8�54f���{����O~G����Yyw�Lf�)	R]��$3��߼�	��>�%r�viՃ���*��$��m]��57s$��®{���\�������N�S#b��T(�@���`x-�Z��l~U�ZMq��~W�w<���/׏ϰF�	"����G#��z��
���Μ�����<������{������-h��~�C!�<�N������!��aë��C���L�\�x�����
^�����{�0�|�wq�
B�*�x`�.�\{+��y�;Z+Z�q�q��̟,��Z8�������D���GW����CH1�?�?�sL�Yh�����	�V����\6�0rv��4�jv���L��ₐG��ݫ/�у��8�B�BŔ[�y�0[�e�`I������o�0#`��n�J/��}��X.M}��ҹ�D~��d�C�4k ���A78������Y4݅r���+bĩ��y����/��DN':i���L�������=�b��~�d���P !-�'㘕�S�@�	<�f�D��A��]���*�|u�`��h�|W(�������B1�/v�����فs^�Z6������g�^���KΗ=sJ��tF��T��T���'Z�v�Kj��_�U>��m.���n�ZZ@�Q�� ���=��\l�4ƅ�w<񇓓���`�<���v�c"�0��>�y���� Ww[���TD���4�]��o��ק�
+$wm�� YB�̽S�6�e����X�q�En�q��c�~�}���3~cC�8E!	�B^TnzD������D�0��[Y~�����<瘪����~���l�6�石T����d⻒4��:\���Jy����xM���c�./��m�2���ȫ�4������m�I۰�?	f������F��l�X��22˦��lo�w/ĝnB�����_=+4��Q�ҫC���R㺪��e�4=�H`��������3ĉ��%���X�Bg\����tƢ٪�h�]u@2.iq�F�}���)dwq&�t��������HI��Ո_�.@�QT���/�L�_.�@sh�e��Ñ/r.��84�FCN�B�����g�K\_�80b��'(��{�P{�e�Qv\�S��\ ��ئ�~�����E�v�*jyl����~�����1�mh��8�Cv5����8GY�O�GEM��Y�����{s(��Դ���<������]7�mAg��lLz0d��@_O�Q�d�A��]Gw�u�Fտ#��w'��}�S]^�!�?���~++��z��:�c5;tm����pR���?����l���۸�~�赙ml F���Ь~)��ɉ85��pq��)n�,ƚ_v�Pvn���.���~|�#R!VBh*��Gǟh*�

k#��U��UԴ��#�6�=�IM���6G?AE[���8˵��׿���V�۲K�(�UK�E�e�0���b���6?9��w;<"H�����'�w�T]��]^h(�i*CBCF�.�Q2�` ����cz%�<\����� �<�S�ߦ2!�ٍ�5�݋�r�+� ���O5�ē�on����j2 ��e�>�)�^Ϟ���BG�[L-Qg���G���;����qO�6������H� �V��f�-�,A�̟!$!\�B|I����C�}���&3��u�
���B'������ڟ9�kf�u_鋜ڵ���1�hO��&�p�^W-[���u��J`��=��_���lz��ly�慷� 3� ���s��Ҍ����_-������v�|��Ww��		�Y)8~�qK ��yU{���i�[f���m����w�љ@Y�W�J��+��sf�f�W;��W���a��{�4�������*7�v�:?M���X�'�Wy��{�X�PO�l5��y�,��X	z��U�'8����D�g/NjD_��B`���^k�F��pp�z�~'�D��0�$V�"�b�J���J�:�5��Uئ�)2�o�mva�o�����R�H�OkUґT�i�%�����A�(��)��M�Lt��x�q�5/V]Ce�I�T-x�,��Y@B-U���0�}Š�I@Up-i��Kl�ܲ�&���D8b�2�߷�z?��uFI�66�;$Il6���r�ZU�KsVz���7qD;�];��������r3�x�G�]O.]?�v�\t�� ��$�"x���s�Ճ��m���I��	�dFz�>^X쌪W_W@7�Ԟ��ѹ*FQ���Kp���\iH�\r�����\[�)OXfn��%͔�⋿������Z�E���tF_�{�U�yV��xdnxB�.��QV�]��H!��5"3�%4��4w# ��Le���W1uT��rP�A�XJ�VQ��������>�hI)	M'd�����؊���t�� >~X��*fMF���)�9+��F�g�Y2Q�b�i���TE��0� �.�֨ji�<�EĈ��3��/W0�.�(ľ5X�U�;y����O��]�FF����o	�����% 鴬LL��Ä �j������n�d*�$�D�*X��ёNH����R�!'+�Xt��)|�:��tc��ǁtM���������t����`N����u�uW��<l�Q�VZMHm�(=иK��(�z���6n�B���T��p�Fk>�T�2�aֈ<r���ߴ��)��@EIW��V�A�Q��?B	񓠦I/�vhB�CaG�О��Y�����s~(���/�� ��V�&��oD�)��c������>�B�eǾC=j�]є���=��� 2\I�O<.Q:,�}��ʻ�r�w\2t[Nfw!U�r�{��.�]^CoT%2B��@rV�"F��%�+�t�̕f	���'�����:���ը�X�ӛ���H,-I7�m�P"[f��{Nk1 ��=B*8mP"�����uwU/�3�.T�%�n|��B��y�Q��!" ��O�O(!'�t�=�R���f�ӡ�k��.rd��e�V�%v٦��?�=>c���(%I_�B$!?�XQ���4�cA"q �#P���A3�G�dǓ?��%���
f����l�~�����!?���$����7��I/Ǭ�s�d���7;;(S�c��o�qN+�$揞l�D@��Z�̔��|闸���k<�פ����s=_� ��#���#p ���2c��9� �J��|0�"L���5|q����]o�F�e����9޿�@�#g�q�ވZ�j�٫E.G������3�<���G��+[@KE��M!Rv�a�\������Š�ֱ���
�)_�x���O#bC]$�r\4P"�Ugm��7����w��Y�-�>!�Bq<Q���*�g&�g/�	�V{0"���-v�3YE�
;ȱ?@�f>�@��kh'�Lgoy =l����T7_���BR�z�dە����Z7�C�X�zQ#&"380}gl<��Ȑ7:#q6��7��D$Q�&eq�9sm%+o!��I�ʗ-��!#�:1��~�[�'D�Lʴz9:������~�B��&:3�;��񞄪{ncJ�iIʗڦ�;����$��]�cv�A�j1��7C�5)C,M;B)�[[�~�5�A�w�H&�C@%�-�~r��x2TUL������vb,G\��8n��ǖ'���-��\Xx�+>WAH�$.�S̽�;+/]@L$���u;]-�9]!R��BJ��h%R>I��wڅ�Z����ϵ`@@���/^�h� Rg���`\w�q#"��$@~9n�H˦��H���s�e[t���4{z4'����d��>�YڛV��}i@�[�P�/@S�c��MU.���g_�w�ϳ�RfZ�'f2����8U� ����R�g�#!_� F���7:��""�w3��E�%�hNPV7�����wT���8�k�e�$�I%������k�<ߒ`�(.��Bqd*-��Sns��ĉ��̕i�[C�@+M-1*���ą#W����383-s�=���������s]�jJ�8�)(ȕ�.m�s=�P���g/�W+�d-�T�L/'�����5 \�|"����f���I&p����*�\BZ_��M����-�8�t�Oh���]���/�Xmu��&=a�[��>D�(���%����n �;�|�� �$� Qj_҇�c��c��G�y�(tƌő}�S��Wb����k{��E[\s���7<2[/̣	GǠ<N�N ��"ʧҢ�ր<8,��BA^-���q
m��񅡑(`V̊���@�8���A	��1�7�sZ��-$C�<�(�{����[i=^�!n8i
_��e��1���kE�Ӳ�s�������7ʯ:�l'|���n]�4-��3,y���7�BDs��Ŝ썙E��ͅ����R�q�W��,N�l�lƌ��AA�d;>S��|�*	C���+�bL^�E=<��2浦�&��ʬ *�$��I����!�= ���W����W���$!��z@ �/J.f�b�9N/���]��۩S�� ɾ�8�/�]���j�ʑ����L:��������f�N[��[���ߧNnI���j+��R4;du>P,0[܃D�hw��}F^���/?5�����t6	p5�Ӿ�L�o��� p�QR��-���[s��x����ˎ�Γ�������G���@gR����'I$d#�q��+�C�@�$A�"��LJ^�s ������u7��9�T�D�M���m�'O,�մrl���q�3x�]$8-�ǋ=��j	��qz��zZ�(mK,���{�r�*6�^��"��C�������I�ܱv����o<���� `߲&[VUs=9���Q�S\�"hRX�9m�\���e ���㝬�+>q��I�����W��穳D�/MyGa�8�Ve���+�5����@�|�Hb��B�ʚ�!��j���� �'D��k/J���mo�J>r �ZM4�˯,�h^��X��j+��*�3	Zr�݆ 7֤]cc�[��]�SP�-��rGz.ۛqN#�>�ַڼ�V�.��y�t���/�������,M���V���.��Sڶ�����D�z�dU���W�� yP�Zo�Ju#��$(�/ո"��E�Q{z�>�O�Ƒ��{5�jJ��)�)Ƭ�5�bDSL�' NP=�k����S�/k� u�-�a?�$�Iw���3�*�!��I�����^]��e/O�re��VGLx]nʴ`�)ʧh;u|M�����'���G��R��0�˲pt�Vy�!�ب�K�j���8Y��E�ڃ&Ƹq�53pV�ct��ܣ_��L��L����<��;���W�vg����a����?/_�=�� ���9��d��8�%A)�o$[㇏Sֲc��~��]1��o��J�� o����d���$
v�Kd��s��[��W�Yվ���qȾtEDŇ>:��{:V�A(;��Q����W�}~rW�n�θWk�@���8v��2�^Km�TT�N�f���"J$Ĥ�����#C㰴[�9�*����n��x���}�.G4ڴt4]2�œ� ,e�s���Do��T��O)��j���!�٬�����(�</��{�g�o6�I��^��]h��X��R���ܻm����91�\D�9���9&�i���G�nn����S�5�(�iuA��r���6��r���HګV�t��o0mc;�v�1�_@�:�Gj���K �@.�պeErjBeڣ(n�¥U�Q<9����X��:�` ���U�J�0�q�:���o�Y(�U�F\�����i� Ֆ���p�~��=�˄��˱�����i���\����F){�k��UG�Hs	2�ZC���u��c�s��,G��H&�tT{��l��HT)�G@p�γY�uU���l�������g�����������f�O��y�R�F������f�튺e$zL��	o[?��7?|�(	�	�IWQ���0"SS�(�Ȯ�"�L��g���t���ȱ}V1�_O,��P%R1�:)�q�8ia6�-��*���#7��?1Άt>�3�5���]���Vf��N73߻�HQ��+3�UVQڟK��GrR5��v�(�^g�׎�1����<K[�WE[���jE�<�MO&�\��\�
~�ϥ�MK�8;��o=|ȓ�<k��A�Wvp�[�p �9DYz���>����g��������1fb�Q �����]��L#A�x������Pi�T�ݙ�B�0�t�;T�WAn�W9�?����+��5�z�Zm�ԡ���	����'�K8�0�����%_l|������i�߶O[���kh�	�f5�O�N֎���a������P�_��T��iqXZ)uTl
A6��ؿ&�&��I�w+��>�ؽJ�|����)(N�=����%�8ջ@�\(��� ��K|T�:*p�-�����؋XD6�^�5/8h���.V�AвX�_�yMĂlu?�R ��❪^�������_Р���4@W�����C���\�h���յW�<%E��S�7WG�����j6����޾���R��P��`|X�OKp�[��n,6�҃Rnl����%��q�{������H�>���$_k��w���-��J]Oԝh[=������~MZYn�Mj��K����`|n������m�t��g����0��رx�v��!ƺ����n|wj���㩡ĝ@� �q�ӛ��Σ�@��d	-Pv���3�Y�vճEܕl�+Q<��6����|���z#G�����&i(,?��b^����ޜU�P�׭	���,H��1Gby�!�Fh�Ccӑ��c�q�qrV�v�R�
?��@*w��f��w�V}��4	��1�-��t/��=�:a��2i��{<��-vvO�+�'̓w���	���VP0���Ρ�С�z��
��s7��n��L׍hy��u3����I"3������!�O�o�8c�+�Dm��JL�>1T����a���*��4��p��}/�v�*�G<7��ǒ�'�t7�6&�ls:�����w��;��7�C� �Q����NO5dj�Ϩ�:e��Z_�2�=��\��8�SH������N>w���j�Yc�&o�$�k��ų�$�;6��	����_��_������7���6���5�)�r�PK   G�rZ�SIM7#  2#  /   images/7346828c-be13-4248-836b-104e84d3cd43.png2#�܉PNG

   IHDR   d   ?   �m`   gAMA  ���a   	pHYs  t  t�fx  "�IDATx��|y��y��u�����ދ��A� �)�$��H�*QDZ�Q%�Vu8����Ju+R(Ub�)Y�eKa�DQ�e���A�)3�x� �� ��k��.�>fg��_��{�u��.v������t�;���}��~��?���q�1����<�[��I�υ����/(�����5=O>q���]�:B�G{\@�WD���PD�k6nC�%��C/`.�@{�)���	�d���1#�LFQd���l�.,�A �B�)���}�6,V�x�����X��}�?ŗn�^��}{���.bOQg�
Q���	�}eiӍ�x��6�K�%�a�4GB������>|�-�FM�𵇿����B��o��\�cۦ+��"��ԁ����Z^ʕ�H��0"&�+܁%��kp>{�j�_��k�eD�	YMt��V�uۥ��%�Pʸj�f���')�C���-����г��⢨��
�<����������FŢ�����K��������5R#��.v����9���ez0�����=�����a�c�0�c���7�G}���>Mt�؇�u������(F'ǈK�h����7�,ɱrC*�t@aaf��֞�hk�����27�c��=$���X�9o�e��F8K-�i8��Kϳ=I�`���a�1�O�}0����yҧ�CC@�kLN;�5~|��>�q����)���1�#(ғ��i���E�+O7�'#�����N v�@�ИO4�0R�ɤ�]L��Y�c��+�*����FD+�G��5���n�9\��TǙ��5>�(����0��Lz+�o�Q%��:'l�rk�!�U��k���G���"
U:��b�<���z�H�|o��[�1��{"��ȫ'��A�c��H#hJ��6Ĉ,C<���_�|lY���0ӭyvcp��F��^�J�͎����Ib�B���#!���D���[E�C��}��^���.#�x�d��`
D�J�H	0N�Tr2!�PAkk9/0�*���F�8%6��(W��m0����2M7�O����_����>V����o��C	��m/19�8_J���,V�\��:SC��g����Il���J��*���Ȋ�����@ԱV�;��؁{�^+�����5���1�_ip��}@����\Y�O����Zq?��g��y�O`E�N��~e~[JZal�� iM-�Y���b�x"���K�ׂ!/g�ę�F9A��w=6�%d_jϧ&¸(�@n4��e2N���ڌ	�\�d��y�Qh�0�B`d����q2�՛��\�W8!Q�rץ u�1�7��lb�	K���A�HM�ܡ;f�&�ط�e�J��b=.s�3���PA�LUL�M���8qnֶ��_�W�d�ږ����^�s�כϑ�"1O��(��kl�f��l��*��e�nb��@��X����y�ú���Rlx��c�@���c7nfe��({^7�7�4L`'��<͐�
�D�L�Ύ���]�:%����м��0D��\8���Ȥ�B�q�@[D�R$���e��C�D��nd]t����h��j�f����uH����BK1����{t��;�s e:q-���Α�d��8��S̤[/8v�����`cZ����Bu�5����[��j�6c���#��p3<��P����$Jwh����n�_�V�&,��!����;�)�����b�W���;��B'<RU%5��lqt��p*9L^em�%�� 4!'1���;!������g�����JDb��b��Ĵ�+K����h�g`��9��W�=O&��@��|�G�~ L�T�V]�F-��g1��O�͍��&e���~(G�;��G`�68ڗh�"����H��Ir�>�Z�6���G��Љ@/�~�ﲾ^/s���w�)Tb������L[�&}�1q�����ƊN�%$�bP�"W�4�@�Xi���c����bso��0!Aaobx8�x�h�N��Ԝ�0F�%�B��n�B�:kcb��%�X/�
T����M痻&6T)啲11~�B�Vb��=��a�P�����d+�&s6���b^�.��lAD���H���-�cbHH�÷�U[ːF�R�-ȑ�T�p����$���8i`m�T��{5�`����!3 �е�ʻ��4�a��)�״嘶�A�t�E�2�j�����x�^A}����JY���bw�>�63���t,���H������r;BO�vj��2M}q\O �m�~c�4���t����DwႵ�h���|i�0O��k��g�H6�Ԓ�,uM(mF%2|�&����^p�.��s7��*����-6�s
��!䱙�����[^8�٦,bq>�m�%�U�;,z�\�3y8��ɞ5�ne�d�cO[�m9�h\69����9��30pL�t�f%�B��-��\W�D�Y{���A^�Y3b{&���j�S�e��L�N�svC��o��J��'�fe��2f~.�N��1�ttz��3�|ǨH`�'�;�f/G�`e�`�
:�]b,�e�a��=GH7q��c�^�ɻT;���g��le��@��[��ש����Jl{f�F�m�g)��֊�pҘ:��� Y���l�5
�X��є:I�Gf�8�in!��w675Y�.@{VM�on1C��\Pvֶ$jl=tJ@w��$N�{69�e�9�� e���2�U֮{fY���f+9 S�@�,+f4.��0c)�L�)`3��<A她,�؅!�jXTc�*����t�3)ʨ�sgQ��G,�Żu��v���k�s��';dM�<R-5����Fd������s��$M~fЧӲ���ό���-�W���&�h8؛0�!}^����tB.�K?�	����#�Lq�Lb�����ā:�����ʱ��7 Nk�H;3�n��}n���9��E� ����<��mtsh2m�=g��I�>G2�H��h<;S��Z���v�za͚m뒃:���v^:P�<%��M�ȝ��hz6~�T㸉��Ʃ4;���v��o�9�)�I���s��Z�)�1�ߦދM�V���)�V�HRKp�������m����8A�������y�,�S���K�8���N$��i���ଲH�� ��Sґ=���@�T�ݺℨJ��J��٦�29.�e�}a+#�e3N?X�~��8��C��Z�8n��^m&J^,��HiE�R �ُ�ܐg	��(�kL����~��f�m�!ʳ׹����h��#1!�0���J���埧�$�U:7)����vj&	R��X!�Z-f[�
ǀ	�4�\M�ws���b��<�u�}� ��!�Nm�g<��<|Ay�d��D崋R��(�	κ��ދ�x��٤�F*��9;��s�M�e��A��Oa�5EJed��iÕ	e=Y����N�%d����JE����x�]h�EPc[0����L)S=B䅿0��C_�=�%��b��ɪɃE��5+�b/�0!}�=nB�	Ӭ�� �f�7��陡R�g�U�i��G�1��{��̞٨<��{�"�7A��ۆV�3}-��3>Dl��2R�P�D�B�pi*��yx�A��r�RT�vO�Qwi��!�Җ��@%��t��u=%� 	��924-;{龋��FK.��ʾC�bf2cqkL-,k<�عr���|k�-y���{3�,�C���I��j7���/k6xdW��Y�� [�A�P��m�(|�$�r��Rg������T������B�Eʍ:D$�qڊ��!Lc�`	����X混±���!5��`*T���a��Z�C$�1�����A�3�e����Ȕq�gÆ$(G���G�Xz]3��x�i��^�����MDBg���e,q]$�V;��9���i�N�Jv#� �8�����H:��P(� )A���992��U�d�n!�?k�
��
�ؤ��(��v6Huގ���~�zk���ҏ*�S1�r��p�臎��!I�n���ƕh�N���fK2�O�4~$I�U���m�����q�`��n��Qvu�]H��8R���h��8����>D�n��6����¢��0ȅ�3�?��!���.�2�BS�������E�:�@�=�����2T��lک��BOYS*	�D}���%e@�z[P?["��盠��~*=\5ρN��T���'���v�cۍ�^2�yT��)Ag^�>���*+p��T��KmA�g'��:I�hg`���U��Ʌ�v�<n���������AWjZ'�q#40D�!]v�\�CX�&��@��'<@��R��Rh��b��� IwD���>#�cJ���$-�Pp��DG0���׭I��� y�����*)��rq jR�ɵ^��$?�)��9��󒚗�1�|��͓�1PQZ����tm�&���-ЭƢ8-J5ĬU�"��a���B0�U)�t���"�j�C�Wz����mY��#'��M[6_���h�����Qjk�ѡA\z�V��=2���ۈ"���c��]�º��>���N�[J����,��+�l���Y�MMb`�%�퇎���ۄ�{_�UjA�?|��~��JAݙ��(����m�f�1�P�%�7c|l=�6ɯ�Q��h���("�v���r�6���N��F񼥈��r]���o����/w?��N�dˀ�A������H�Hs��/Q����!�����䤫�� '�FѢ[����pXs���8=v�a�qt5�lXA+�@���T�Vހ���h��	ynm[�sg��l��Ù�f�*��ڋ��I,���=��V1Gsmq-:Z6b�~�D��ĉ� �aWl��禠j��nƾ�,F���Mߌ��	�����\7����&XH��ҵ�]*�U|�N��*�Cr���������>R��J��ă�4u���VR�:CN����.��T�L�*s���ƾc�c����7_z=�я�R�{׾?nm����� ~q��x1�'nx/�΍���I��7��-��o_s+�^�#3�q͆���7���ɰ��\�N�?X��#��S׽�Ƈ0�8�ۯ}�H��fO�o�ֵn������߀��^C5�ׯ��y��1�g�����១�+�S����\�^�41��O����f�A��G�l>	�<~�m���[�1
�A����7&�P*��N6��:�%b�/Ť�æ�Z���IZ��2⭓��e�n�Q�2��:K2����Ѧ:�_�C��PT-�i�E��<:U	}�n�:��]hG��z�ݭE����Ȅ䱦��L�r@Et�!WU(�E�m�A�ݥ��[�Fg[ڋ�(�Zֵt��ԁn2�ݝ=�G7zs�OWִ�G[ЅK��1�O�ף~����~�W+�ќ��2/��;ߊ���ˉc��	�\�\k 6#��1�`ϣ�,t��$�{���Է��MW���#U�?҆I*CP����g�2;Ӊ#��!��ƃ��5y��:�|Eo�\�t]wW
��+9Ϯ�N��̫<:���3����2��a�P$���N�2�������2�=�ȏ�|[�����&)n'?�$��N����AZ�h����%��]W7 -���dZ[&�z��0M揝{�������/�LtRN������J����͞�H�r$+� c�'�����]��q)o7�,����-�4O�:���lBG���b0c�bX�f��TۢXe����M�7�Ȳpq����ZC���<�����O]W)��!$�3U1[�9E�Z��
���LA�:Y�Q댆�{]���l>��Y:W#�����İ:����W���vQK�w�� ����ja��	u8.���)	uE�_�~�ZE `���K�1.�I� G?7q_��/ʺcB���v?���4�k٤�<�3fFi���J�����X���D^�ƶ��,�3�*��̀�2���ǽw�]�(NM�#��}�O�7N��&�;���睘���i�wO��K���^�7y:H����)|�����A�b��'������2�v��IB\�����܍��9�P�}S���Ç���]���B[���cg��c�ͼ����V���0_�G�����~s�c����~�fgprjc��ZT��+/�_���+��W�pʹ��޸~;~�[�2���~W�-(t��?���	e#GG亾5�x��o�����o��-��k���|O���%B]�"����4{��G�m!j��b�F�
��!$6��I���U��z-.��c��G��oLM4�v��>�S����Sd�M�xqe2��u�=��|v��F��Kn+[��Pr�F�F�8��l�+o��y^��S�"i���Ce�b4�$'�����#���ő#�%�v�(����������<�����/�m��T�̾�,�SĠv����m'l�7���̚�0L�;�
s�<��ӷ�R	�c�S|�)���sݛ%�R�,)s�L$���9�,��/����ö+�Ň˾�;~�V\v�&<s�Y
y[�kC����l���Ĩl�)�:�ǫ����x������1=5e�|!�]�ش�r�R��oG�l�4��m����-������$fqD>33���0����i�eӳ3����]�1�d�	|)1�Tj�Su��sYC&~e���K(�5��|_���^tt���졵-`�̨��|p�mۆ���hm-�� �
����f��Ds���f)�]����q��?��	2�����}�:Ic7E����p����]��%B=���o�^y�6<p��"���/a��>48��7�[_�:\��ib⌤{8Z�ב�G�DI���٭�*1�^�lU��i�̤�[�Gh�'1Ec-�^��g��)c��2FGϒ�����C��䌘;^�J5�A����Պ�������,F���Tq��w��dls�fHc��C�:�^�g?�Y����������������5�{�"�:/���'����YT(@,�9�!{��� ��$o�菴�^�JZ�&m��Y�Zze�SU�h�S�vZ
o��	��j����k��+�`���d.'H�*��?��ش�2<�{��Ǯ�؅
����r�I
�<�'�fh��M�=!o>�S3F̒�E�질A��څ��)��;TX.����?R,��C?�T���I2s�"�sm����!喝W���J6����u"�N��ˈ�� )D�[���&��ȉ����C�g��s���¡CE�����|Zo��\q� [�
���u���9w���!4�+yu��%�쥀��n������'��C;i�U�9L����=x��#�����zA�=� ۷o��?{ǎ��>�Z~��w��w�8?ɚ�L��e$�mS1ij><�b�����t�5��L�����g��0EKK^�NBu<��O��K����?�"A����۫�5��X��/�]�Ǐm`Iq�yb=�쳂�����Gk:���}�z׻�[��/p�]�Ė�[����Ǐa�M���;q���;E�(�8�p�E� &���BƼlL����uE"����j%������P�ț"p�ǦH����K6�된���iXM��M�`�Ԛy�%y��f�S��+i���	���_b���&��ƶvϞ=���?N�B̩�H_��[(z_��}���~{�\<p���ǁ�ϑ�"r�$���)2���8}&B��D�HY���	��bq�|	�SSY���ɕ���&�G(�3P5���bf�B�N�y�^:�^�֠��'� q�xǭ�C6aﾽ�hD'[��z��0e���תq������K��]��1'�&Λ��/7`S�A恃���A+�*�L��5qݺ���$ݓ<���H��	� TȄ�esI������}r_��
�y[{�}�:@gG�z���8����+��9�ܹ[�n�W��U��y���:'��5�a��:�Il�an\���\���r�|筸����;��_5��'>��_8Hq�:|�ӟ�]��v?��H�(Fn��W'{��h`���q�|�~tX� ��������dQ�D�Rj!�kbL�$s^�T�r?�96U�7oF__ߊ�^>�/�9��j�1�������(��'?�	�x�	��h�̙38q�8-~�P�9|�S���3�����à`����0۠(���ld
�X�8�/���cϓ����/�<=�7]{-���L�7G�88���ߏ��LLN�Z�#/��y�x�b��:�K��;-!��E���!~~�L��؁sT�Rh�8��o����ѣ����9��/�ɷ���2����02r:q�|��?�e
�q����AP� �On���� ��<n��9*H��ٻw� ��c�P'�Oξ"�L�m�k7�P���B��F��
7���m�')�;;;+Ro�I}0����;8:fĎ��&F�8�H,���a��q$�����Y����W%���ݻ��(.����@RrD�Yxx܇�0�yӵPL�|K�f�da��xq��.9ϒΎ������W�����o��>����[n��o|C���;�i�1���o|���o[$���n�W���w5ͅ|A�'�|Rb��|�#�ַ��믿^b�{��.eM��c�waa!�Q+5W3�l�GÂ��o�-Fg����2I��}
�h�N6Yl*X���LLL��oF]��9��uS�ٿ0 `-c�߱c����C�8qB�a�]�efʁp�*�lk`�rA�k�����|=3����/�T�r4)�~�G�裏J�������h�Ì� ����7ΞK����Z�a�\�ǜ�e-a���#;�ٙ�$Cސ�UH6�Vk�Q��ӳ	�r    IEND�B`�PK   ��rZ�c^��  �  /   images/7daa3674-301d-466b-aa13-7b9309bd01d6.png�B�PNG

   IHDR   d   s   n1�w   	pHYs )� )�;d��   tEXtSoftware www.inkscape.org��<  JIDATx��]\�U�����@43\�����
�����̑[��Ie��ܳ4g����L-7KeȺ졌��x	p^.W���z��}��=���s��ʨ�QXX���/����'R��p:s�M�>��ܹS�Oip+�V�۷o7���w���S�R�fef�����?x�@���@\���z����}�:��z�rC�8SS�++�6ttr�Ӣ�֭��x�bj׮9::R�^�i߾}Dj�OM�F���),(���X���k�(.>N���ѡ�ݻw=gϚ�9s��|�]RR�~ZZegg@���ED�<C�;T�����JCC�D:::dhhHfffLF������ٝb2N�A��\�Іf��(6&��RS�b�J:D�biﾽ���+����hݺu�y��}�֭�111���T����|1r�pGW�7����ĒE��M��M����]�6�I	nӺ�a[[۽|��={��0�L[�)5J!���'�#�Q�t��	;g��~~~��z���q:�L1͓���RƒB)))����q��U�#G���ܹ�M�^mӦ�6s�;xv�\�n9�8Ӄ�D[�!5�J��z�n�N���x���G>�ƍ�/(8�099Y��Q�(��ZZZ������B��}���{�� �={��`������=y14$�\\](�A�hguSm= 2�̝C�ƍ��={�_��r����F�ٗ/\#++��I(ؓ�Djkk�����1P�h�O�>mx�ҥ�G��R������������߿D�U�hlBb��
\����ݤ��fy�=�z�uYNN��pt��!�?���I___87n�@IOOO�����`ǂ4BBB�:y���ɓ7XXZ,hаA�-�^�����Q(!������h�z3�f�'M�4�ܹs��5E�C�,(�	o
��i�_��xݤI�;w.-[����&�fY��Q|}�����;v
,�,�5�k�+�m
!�.#=C�������ŝ/��C�u���V"JC��z��	r�߿O���4t�P���o���Ӈ���͛7���	;v̔%ƿ[�n�Ə?v���Wq�i�id`h�o�	��
	!�D�.��0���Wl3ta�U����@�ڑ ���_d ����t�R�ѣ͞=[H>T.���>|�T��ﳳ�E(¶<!h��ի�7� mm�m[��X�`���b+/���$@�M�2EHΈ#J��ԩu��QH��_-���]~^��܎�݇]�4�ų�ReB${q,�\B�%K���o߾���*-OTp7�5��H�۷��/ )�+W���n��'�����ɳؕ*U�޾};q��a���;9���hS��h@20����hƌt��)��㏩E�%��@�AEϛ7O�cǎߜ�5s� ���|ҐU^CT��@"�U�VQ�={~:��O�<��$�6�g��1�@��������ԵkW��,--KΛ0a� �G����{���O��j�_>���J�T�IM�\����ӭ߼����|^U�� %,%��ޢa#J�W�^�ꫯҘ1c�&{k�fL�1p劕�||}*��*L�d��n�
��5����Ґ��$ =߼ys;vl�s�☏��޽�Ο?����E�gϚݟ���CW��W�|!��ѣG��G�ӦO��E'�4������Ed�8�<V�X!�d��'q ���_����w;z��K��V����/�~�:q0D��4n<mڴ�l�t^2 ɮ888ЦM����^�� i۶m��w�^:q��B��LLG&3}XR�J�mY}}㯾��'��,���B�(�������I���A�v�Z�������f�f;�|:�CFzF
��ix"!�`����M�����f҄��
)�G�#�^PmFFF4�|ڷ�������: }�4�뱄H����t�̙I�.�/%_f�S���R�q"X,�����B�8p�v���}�d�,-OT]��ݘ��~�:5ukڊ�⢨;Q�2ٍ'�ԩSG�Z|}}���@�*偈��?�����=���`[�����Qx$!R���H����.ԩ%�,$R0<~�xLj��K.��q������'z���O"�DU-^L��z�ÿ���jQ �ᨨ(Z�|���1x�`:{�,���O0�-_i9����I�G���A
6̮���#-P+�+��׬YC��Wy,Y�D,u
�={�����o~4pP��<��0=��3���2�/��0`�A����N �����`�֭�2��R#	ez������w�� ,D����RWv�����pvv����~������挋�K��J����p�גQ	�[[[���/ń����C����_����ܶ}یѣG�������B�a~����V]U�POH��d =u�T��������v��i,�� z��t�[�n�V-�����˗�����{�s�C^�ĉ�k��	#F�8]ZJ�z����~���?�[R���t����HB>����[$ 9z���Dߍ����`f�R�͇���j�JG�!M�^�x�`�7n��9�۷s+���Ρ_�t��,OOOqL&��o���6�IK*kQuHű��,�v{��O?�s�Ͻ7w�܅�V�=��y�gSϓ����[��#f���t���9�{����޸�����#�y0!,�-���w��v�yI��l�)�a3E�O5�
��\������9�����>}�t�_�rK�d0�[�lљ���.X����J"B�N�{�ZZE�jE���]��NɃ���u�x�&�A;1'�Pbǎ�����9xǮ]�օ��a.�e����]�[ᷜH�!M���446"==A���t>?����Ρ��4JKI�L�ZL��]�D�
���mۊ�F���NY�Y�"""��0)����:�����paz�d�zYO__�KOM���22ҹ��s4��utuɈ	321!K�dbnF)ؤ��$$F�҂6a���͛"�ׯ_���@Թsg�R��_g_���l��1����=����nyH��Eݺdja.^G߹Cw��!b%N��-6�}F[G�,�Z�m�damM�L����l�J�����4k�L,��y�f�1c�,���9�wÒHU�������̄UO*�
�d� �=I�ssr(2�6��Ē��� ��}C�a2�32�F�� � |i Ղ4UdT$�+�VW6�b�(��g�d�R������>w�z�*>�`�C�Rfz�4iL�Xg߽!S�F��BLR���1�����J���dmURW�l�M,,Ȅ�Ƥ��v���ԫ`�Ԋ�����[S��zt7"R��2 m�;y�$���P�F�J��M��>�@'(0��,**�	쇪,�sլ�ͭ,);+��X���>\���H���ۓ)�ĸ{JS]R�#�@@(A��������%��� �Sh`eef*���5޾Ff��
�(U�"T�2��;�����E�i���.Ā���.2�\n��
�����p@��!.&�48�q�|wYR\�6�Lҽ���j8v�!:���#ޓb(8U����E�JeV� ���o/�]T4R��z��NBCGd�9>),�~�&�w�ok�$BDa*� p!���2VV��
���z���DR���+���C*K�;H�(����]�z��=i�#�eee�rssuIE�ѫUG[tv�V�*�ŧ��r�X���e�7��B"�R����	\���i���H�$
33�KZ��
�	��5�2�J�#P�X̓u� D*���Z���0EP/v��aU���EG`*�
CE���!�^z��/u�MhWͻX$RQE)%��Ջ�)[;Hv�����ui�j{1�H�jhTAA���ji��R]�U�^k��K�e ���Xك�]�T�p!�����7j� L(���S����%tj���c0����Ҷ\�t�u��oCR ��t���rp��)8�55���XD��s�+=(����`.
˭�|�����%�zP�l/��efiAV�����>S�c	IM���lB��+$1"������(��pW�W�t2�D����RH	�u�O07
���	H;����M@
s-333���J�j�����ř�������kk���--)eg����f�i�f,��Bfmm7�F)oT��y�G�p,NH��kie%rN�7Þ9����А�7� �X������}��Dl�ƵAb�����K���qall�2�H[qGԤ
�o��Ƒ��69��_�NDdI��� i�֢�ȸ�EGS���� %O�����& �-�9���`Krk�tx@qw�R�vԨiSֳ�q�VI5�� �+��ͩq37���R)I�5N���0�H�S������A�96(�?Ɔ��mM���gR4K��m}�g213LX���EIjʔG �˖mQ}V 1!&��T�V�����ѲF~P�N�w.0�ŚS��I;"���;�#Ȝը1��+��<9Y�Ę�3RP���.F@�o�O��bˁ�a�D��.u�f�����m
2��^dgk�gÆ�a	��������`)dM���@̩�ݽ+�TH����PCP_пy�5�%B8��1D���F3q�j�?�M>n����*GY�W[����_�5J;��!�/Uٵk� �PE� +#C<�h�KI���\�9�81��_���Ey�B�T� ��@�q�xΦ�ɘ4��ҥK/���.\u:�l�"��H��)�ԩ�9�b�n�Z�6D,�-vً�qL]�� ����z��6{b�����>GG�ΨH����w�+�TU�PD��#^�)̣��2$uղe˽�7mo�~���z��AOO��7lؠ�ſ(����N���q�*��k,�^�p���k��	PE�8b_�zu�/����O���8?��#��P5Iy��עE� ���ev�BT�;F��m�{xx�D�ˇ~H{����%Dq�t mҩS���{p B *(�8Զm�&�bl(A9;,��-�P�^Q�K�9���9 �ݯ��J����!~��@A�VG�l�s�t�j����{��E��L$T݄��(��-��K<Liu�"!�Fa�X�a��� ���Q+���ǡ
����v�:y���Q�`ذa�.9(�����И��pq�U�(��T��@]�j��n�6b�-�C$�)ٷwE�D'���{ف��DG���H�F�mHLU�d<d �1�T����L���;�X����ԧ^��-�Yf�*l���+������>��3��o���Ġ����6��9s�C]�k�.��W�zC�y�2�@J�\��������]���?�]? ����w
��$�"�,����~}��߻wo���ʙ�9�M�Q��a@�Ã���@�-�CMA�e��EJ^V�����Ǚ����e�)��D�,�`����|���lе���ؒ#G���)�"�Z<��lӦ�����N�ܥ3��S��������1͞5�����°��y�Ӏr��ׯ�lP���jIy:�U�Ư��^g͚u�6�1]�HB�;��_0/w�w�^��Q[U@JӦMkIy�B��z�:�f�7�C,�x\���nL��b������q��Ӊ'�ɫ_�Ư�J���j-!�y׮]�YU�bg)OWG��Z�}��O��,/�N�N7|}}G�]�u��I�3g��}�� 60���C_�.��f�4n�����q3�&M�4���y"!"\\�������޳�)�Xǅ��K�.��*�n��`P�� �Q�yx�(q�RUUS�	:��=z�,V��q�i؍g�� +�׮[�N����?��aRǈbQ ) J���TLyR$}��Xn��j�HkT�� O#G�\��>�;M�����B�Md�2q{���ddf��+�/�i����X��Iy��HE�UR��� �>|o�~}}��3���Q�6T�ɋ����6l� f|�ƍ����	�`V�I��q�ʅ> H�6������|h�F�.�#�������~���;6n��s%PaR&�et���0��#F�x��"�Ҡa�J�_*U�It4�����.��/��6nO��e#���6c��^��H�x���D��+��t�,�y�"M�5��z9|�p��5k�����I��, �.���[�N�w>0`�pX��W�&�U�X��Q��`��ܺu�S>�b�ᙳg�ZUu���aR�վ}�_��}��Y#�$)�l��T9K\�r�Ad��077�w>4�������KG��֋Z�R���n�L�:uk�saaa���C�����\ӯX��GD��+f����?��		Q����fMY+P�:���<�s H:�:���*�(��>�~�j�ՙ�W�.������ǝ��pL�9YQX"�+��:t�@F�F��y�B1���7�/ER�VA233e�6o:8gΜV�yL����	�.]ҕ
5?/�HD }���!o޼yBxx�KPp��Np����+�z��)�\��G���bŊ�[6o��G�^AAA��U����ܛ��w��駡C�Ng����fWgm�j��F���ү)*2*���gz�͛7O:u�T?�/u`��V�U��}�1�Q�F�����������?����Y݃�Z����+R�HD���gҤI�����ݳ���_g�m0]���Х�ɑH�G�rIM�4�n۶�O}��Ycllܦu���G�����ɒ~1N�N��GEE�:}�%K��]�r�ۙ3g��]����۷���G��%�A�K1�X�����Oe��D�v�7w?4y��W_}U���)Vn*�STZ)k�R��l���ע��Rbbc�������۰��x��n�>��u�a|B��ւI�U�o�|T�_z.}o�b#,�v��mmm#����jѢš�-[�s��zHLQ��h�� M��eA��Kw F�[]��&O�G���n�~���p+����s�εd�i�4!>��<En�����Տ 	j���E#^]M]�I��[Y`���� ���D&!��u�@��c��!Ӹ�^S
�7�m���i�%A��SeP���K_4TZ��ݩ{���lv/�DGG_�����9�B���i��i�V���\.7���4B�BV+"%���������Ke���������D�Ç��{`! 11t�ʕ�;�T *S}���6�ɉ��O6l���$d��di�:�B��\����i,c��u�3�h��#ϣOU�2��GE:�qi~5��#�|T����y����&�ED-!*�ZBT���j	Q1��b�%D�PK������Q���~��"�|M�Dz�P��oL�C��[�"����~��8�"���ѝo�c#?�)��L�c)p�I    IEND�B`�PK   �rZ��p� �� /   images/7e81f6ad-0912-4ff6-bfc6-e58bb7840941.png�wT���6�qPDG����>� J�@��R�FjpP�A@����& ��&���"=@BB�{��=��������z�g�������>{_��{�s􅞎������@ �ݾ��>���`�t�����1"���mã�8z�9���>�e�@�|�9T��� ����������B��=tu�yd���!��p�8��������_���/"_�c�?Ə�c�?Ə�c�?Ə�c�?���#x��ap3 q�1tS����1~����1~����1~����1~��+���������f~��ռ�䣊ʷ���������N��W�e9��;��Z�����=�����/�̍.����;��'��Xb������jR��Rӭ7�_��tg�WQ��;G�v77�Ҩ#�S�v�P��d�^uw���wE~����1~����1�?��C�qLw��J/i`���[1U��*����hqE��R)Va��jt˗/�,vLe����|�)��*�N}_CW~�����C6om�Iu��Fo]���O���j����Ӄ�adF�� ɜ�)jϣ]�x�A+�n�iz�����T�'3�Ԑ\�c�t5��^�ih�_͔;�o`��&����Y�O������HA2������h�bw�χ��k�N�>aS�淟�~B�Du����X�<�a+l#Z�V��yf�._{|og#����n��Q����:Í[�(1�u����I���7�<�Η}繻���_��ƿ�lB��Qx�ING�^�Q:�`ݦfB���úL�?b>߉g
gVO���$���d�W5�p��s=�[�-��d�z%��`�zd�����S�
�2NU���go���3~ϋ=��#��y�-�-� ߹.�2[��.�u,goz�&
rZ�T��88���<��Z#h_���İ���uX/�sTF�lG�h�[��t�ڈ�i<��3\����e��o0��p{�R���O|��b����t�� Tw���|�e� �')�^��1�"�c�Y<�-a3�ç�fV��A�E@Z^�S^�Aś����-�_�b���a�C�䩡���&�@S=��R`�/n7u*�K�f2����z�̂*UR�Xw����;J���mIW������Nz��p�l�;TmV��Hi��&f�ee�RX�_צx[��6&��4�7k=�k
�P��ah�c�{�h��rvv�����ͩV�K�Ֆ1;W�g���s:�8=oQ>~ؽ�|��["y�8�d��9V���m�T�Y҂�_C0߮mH$�;.J��s'����X�Էe�:Nڥ��R1�?�dV���+'����pזA�G=���3��NP�jc:�����f,� ȳg:<k�\Vj���U�b��h�zE���n�(Ѱ?%eHm$��:i��QyuYK�������hs[�9�v�E�}#��=AYɚͷ�����j6��~����×�j9������%�I�±��Ð�m_X3��٥x�6�4�� �1}*u�:6[ĺ|�i�CI�{K�\��-�ӰO�� }�/}D���d1�6�Ű�Z[��
�}G�2OUg�@�\��n䊳IKA����	��~y��]��>��\7�(�qj�?ޛ&YX���Yf��קּw�r�e*�)��Z��(
|�KI<񓳨�r@]u��5o��
vL_d<�dL�U�և��R����T��@���_��}橒�b::c'h�m%`��t#߿��B2"�'�%��+'���g�ZT�+\�y"j����կ^�ʙ�P����#��{�ld�p1�y�?3��˫.���^+�Zm���u`�a�Z�]��-��]��PA�9�}�z��k��o��ru����i�&=����/(��}���!O�Z	�gg��oQ�7�	�������n#�~1��|ʘ����~7�����V���Ɗ��<yD^��bd=d'�S�$�^L{�ؖ'��1I�v��˯��uYW���Gf�U0"�뱱�u�2�ל�����5��
����j%�7TKj����6+k#��'��{L[~�l�5��	��I��gU;u�,��r�{ ~ G]��$+(Ĕ1�VQW瘋�r5sp�tv�:���n��������%����0�)w9ח�rRRO'�\�|Z�A Ѷ���S1�ڔ��	�@�־Ɉ\]�tV���6��U>�WxG��n�>D�J�9�ݯ &UlX�Ƒd�p�v�a;Vb|�l9aX?,�y =�9\��yI�/��|���Y{ٹK�"��Dٲd>e��k=M2(�R)	�t����A��|��A��msKd�zr�V�@Gk�
�ѐb��m{:q"��s��C�SY�n�U��`aف1ȇ<����Te?K��M�;��Z:�^&��G�/mΑ�s�ܻV�h��{x�}���;�Z�B�~K��ʻ��	)i�������d���:o�~6������s���
���((P�n���ӂ�ac���l`>{�8R��l���+buڶ�j�V�4���9�,�ys�ҋ �R�ᇠQ�.��m��~���ѥ�KYLO �E�<ǧ�RjG��د�_iV���:F��u�[mqkG��N��y�ٷ���	���>~�b�IDW%�*a�$�]<�Iſ"�D\��5m��F̺���n�u�S�I�,�c�U�B?iɇ�	_�'Xơ�O�8Bmx�̧�u�֫��<e[�\��b���|���{�}���>�Xn���E;�Z9&�,͉Ц��]�m�������a�7�خ	�l�"�u��YsHQ'�{g��=��ItouRz��ϝ>��1Tc?d]���zJ�LE�C�}p���X�1�I��.I�J��55Ͱ�lw0�X�Ī��n(RSC��=Y;��ۙ�S�A�C'V��Hl;u�PT%v��١E+X�6�F�H vt���h�I�M\I�&!��/4]ޚ#w��.+2h�(����CV�.�8����s'�k�IY����� `�b�K�)V���UϧJ��_��x �=h�c��&BOqw¶�w��
_!ƨ\����i�X�>�ғ�+�u�׊�wO�y��S~�B��ߦy�9�yI�.�*� ~�x[�(M�����3�����ÿ�󒵔(s���my>��7�C��� vx����բH@ɋ�Q�w�)� ��A��}�Fw�b�+����U�^`au����9GR򘲴K���ŊJ��n��.x6j�����j�s+�g�So\��e��Y�3~S���1+$��j]�����&{hnTM��=��B幖ۗ�k� ���џ=�+�26����2�.�
;�d�S��(a����3���#:�;�K�wJ���Lŕ���Z(�w��Xѕ��a`ZBy&8�v/zB�j��"�i�ig�� �����.��w�eZ33�)hb��< QIi�P49�]<Cq�,��,���x��@�>qJ1�g/�,��zѿ��@奧P�N��*�_Э���ج{m��:H&T�����I2�߾�S=a.�p�tX���S}�]d|�д��P�su�Ǝ?���*({&�w���l�ZHClP��1�S�tMzlMdi6���k��3>��T��Qo�^�D�1��ޠ�~K��]V�w!ҖK�j-ۃ��Ui�뽷��W��_���X�9��0w_��Si���.�s`��Dn]����y�7]̑	��E����
U��>@��9|��7�	��k��s�u����RJ�3> I9;��nށ��0%Y��卤)u���Q]�ޖ�eđ�߳|���bg+��v�O�欪��9�2�� 8��f6!i��}�	���~���VC5U�0T�����+�*t���@�K:xM�bt��ux�lܗ�&BX�ˡ�i�������Hߩ�#�0�FE@vt�:c�dlz��$c�k��2����0��B�m[��:Qy�Hb���V�$�оN��jc�_�0��CB(;~Y�4@��^��ި����>%�S����s��2�ǯ�D!vv��ؐ�1Z^*�!���]�o���z.������M�f>��琾�`x6���o1&�-�;|����?o8r��x2<�c�Y>�9��a��q��T�O�jX������38-�tN�~5M����2O�}�ub��ޖ�0+�����m�uv�l���1��]sT���APH�� d3�D�dQ��^��%g�>e�x"�)�r�b�H�
Y#�"iqYvu��|�����FZ�U\�!=�/`F<��v57/��2�g]��������z��+��&].�p�4e>\�L��`y7��[�!$�,f�k�}=�Ņd=HM9�F��+6��hU��T���A���+���..�����Ld�CjJ����m��Qƿd��2��avj���t|��������XGd��"�[�FN����ؼF6����@�g8$�)��2�����fKU���A�)��q�����$��,�iO@��]��L�\>k�V�Q_t���6d��F~�O��S9�K���& �AR˃�"��S����1�!��S+
v��������6��23|�{Qt�!E�eN������
�{�� �dJ+pȼ
ӛ�������3(?�V^c��s�����n��B`�u��7~S%�Kا�A�+����pp�~[���ԶV�9�~-���
���t�2	��VX�g(�R�M"�?�	@�uGJwK��O��X��YڭU�C �VС0lȖ�B��V�N�f���5�����N�Eë�﯌����������$Ɲ�����
.����^�ŏ�{���I��״e_L���;����Q,�,����8���!��Rkq����Ҫ����m�r���]i/�?C� ���"�x�
�8:ٰ!�!��r� ��_̻��ϊ�cx��)�X���D)�� s�4�X����}�Av��,з��"�7��{�P�oU&�o� ��RQ���|e��\Eo�N#2ԑt��/fӟSJЯb{�¤,�C9p���A|ښ�Q�.U@�;��>�ttl�V"�#6�!%.8-V��@��@��W�����E�V�UM%�Hn3,/=.t�!�����!P��W)C��֍�,p0�b.#��U�l�Ыk}mTz�87�6!�������W���F��BWͅ�r�4��[��Z�sdF�V���IB?�c��`��/��1,WD��')�o���x��7��J�6�;�n%��������!c�5�\�ñ���}<�W�yI"�*B��}����,pl��Ímd�C�S�컶H��z��tG���\��T{`a����ۈ�Pes�i]fS�;Yp���-�/�/~�V��!0Rj�=]P��ҏ�=�|���+B�#��6�s���������/�aH�'ݴ3��@'O	1�\_WV��Em���0�����<���òx6����U��l.���&@�,<�a���=\�Ɇ�	�W�h�&s�@�ջG�#�yow%rE�	']1������E���^q�O	�r-\�;�?��4�� �'��>	F1� �ʓ����jf�9�Ĉ�&G@�Gj��KY��tub��J�N&.��#B��Y��铥fÉ�Tܕ7%Ѡ~ַ�r�9w{�7:�=��Da�WC����[vh۩*�����=����l��V���LʴC-M���xQ�Vj�}M�<�&�C��}�='�KB���q�5[je"F��T=1�ҥ$A��D�߆�6@A1������F�{%2���3j�u�E�Zˊ7��2*�g�v;)_��i�rR�R���R��/�]n=�C+ԖWynU��Q��H����>�=�S)(�ڏ��r������I,���&�(ut������I���q<�Pr�*ЭY�մm?��t�����&�߻�E<j�/�8�o s@[�_D���Ed�����)9\�B?D��V�G�����YU��������%�{�-�R���&��A^�"�-�����X�����5�L0���/@Wh�����T�c�mϰ�+4#�U�����x�`�+���6zH��yaڃ�ZL��%o�<G�;]�?Qam�vg9)�̩��΢�r3��؏0x^���'`�2t���.� �*э�qz^:K,��T�z��	R^��{��oE��}R)eʎ���lL�Z��}��Z�Av�m��^z�,hH�w�]~jv�n��7�TTu㴙�֍5����?�:@&k
$*�#`K[�E�]����H(��@#�J�b#JDNя��8oI���2Y5q�!I�w-�ha�ns�2`N��������Kc2%�p�=Z;��R�\/%E���F��G8�&<'5_�%�ғ1�u76e�� d�!�	3��ų���"Z��X2��`�wfIW� 
Yv�,�
�^���b��X�%-Eos�U�ӹ�vބ��I�A����c Z�?��/��R�7Ǩ���]u����G;J\"�q��_���zǥ����t�2�M�����j�hw�Z��"W%�j�d�L�)��q#�*���gA[��J&ٜ���J�6�W�d@�g'|ͮH�\�{BnC9	��_.�,6�^;��?��Y(	����+U���ŻX{�=ڐq��.�䲷�x.�k�JGb� ���rK�A7ܥ��}�+�� ����#2��������Ak�vf[$q9%�<A�b\:�"<e5���J�������$�(��B�X��Z�JĖ49� �ڃ8�!O��ϵ�&FIb0�-���[�<��n�U�)����y�y"������l[KNEgF>���@t��eT��0n~�����Ģ�zg`KE�@�� ����z�l��o/���=:���4?��Q��st;����m_t���n�/�yP�2���/�o]+�dg�\��X��;�>��$�,��$q9�f�ʩ�R�oA��>�����}�Cg3�0k4r;W���W�T�<!` �r;hv������SP�́p���:��Hն���H�Qg��0���M +n��4w���E>����~i)�(l���T����ڻ�q�M��<����oOOeAC�W��f�)j.Y���b�{��y����<7��6.Wák]b>����of��)����Fa�Q�qګo^�T�JӁ�A�'NT�&���T�"O/hᜧJ��襕���y
B�Z�:$�\F�s�7L�&lϋg�󅹦�؀�v'Tv'��ن��a�@�$���q#S|üDx	R�z�Hp�ޅ`%�?q��_,�!����F|�*�����9F0Mw����u�u�w�Ƶ>��	l���D����}�e�n;�I�*������?IN59`R'(QE�����5J�<۪�^����DHJKF�v�[S}o�t`�#��|,7��k.S!�A�$�u����E�|E�Uȶo �b�26/u�
�[�P�tu��]} �3��;�	�}������+��q�eؼ����������9`K�H�99	BQ�a����rZ��E�FN�US'�)�t�s��GYHZ��j�@Ep8�m�n�{���C~�ӭ6�~C�v�I���T�
3)�4��s��%����[���^� i=lS�9��S�
���o�װ�@���X���Mf�Ʀ��O�����[w�N�v|�ڊj���#8�d�!k%$a}�6�;�i�,i�!C֭���X���� {�Ta��7˾�$?����W�R��AΕ���ef���H`06C��>�bn�"�<q�%�1�p�bDX�\�Ɏ��8���W�P��<�|�/�Z7���ą �����>��}��4��!����P������o��	F��Mw��uu��X,�88�5�i޾�cfIs�"-x@`07�T��Z�G�� �#���~�m_��T^b���Rg��_Cs��m�A�f(��继G�*Ქ��{�w~� k���M�̆ {D�KY��+�L����'9Ze%�#�ۯ������%֞��|�4IH�G�@��y~\⎛4����mp�r&vGƫ!,���"^r�
�f�դ����Y���(M(&Vo�ncL�Ғ�~i}�Т�*�ۃ�J3rW�P�+���\�����|v)pU�r�"��s����7m�w�H��y�<�Nvn.���*�;���y5W+�e�x:4KH胝�p��8.b�����jJ�s1�JNn�	��~r#x���_��Ax	�o��[�$���b�nDM֢��9�%��3[AU6l|�B�{�}T��Tx)�N�*�@\s��U`~���a �����I׈�h���c�0�YS��o~������?��|J�����^�n��T@��ϪO�
4���g���|�~ڢ��q���@^]�!�P���`+R:e�K!�?�5���E��xuQ� ��*�!��] (pi�t,�֤�4& ��zk��]Bw�R2���X�c��jlbo�ѿ˿�r����SDt�il��Y�t�N+��59e0�1^;��}>\J#O���p�a�Uk����CV�G��ҊP�:K/��e����P+�*ׄ������ֲ^�aֺ�7�6�GŌab�0Ъ�̽�>��2�	����z�+\'.���Ź,A���IaR�G(X|�2(��٫�������7�r�K��6�-��갲m}�c�g��oħ��A�Z��ՂD��^��j�`#ζ F~�_��b�@��k�	���~Nש���Pi��8�+��ey����@�.��0V޵�oJĥ����� 2�c���	4�E�����Qq�SdQHOF����r����T!��9ed�`��4��,�BS9X(�۲�Ŧ�^��Mr�8��{.�\3�š�M��=Q�[����ZCZ.|r�-�=�3a�+�
$���$�g���B��Z�x�@��y����<k͙/|ỿ�����W>��"/�u:W=K@��Hm�8��e��x�U�-lL�LL�KU�0�I�,Ts ʛ���)�����_�X��=n���`E������s����������s7��K �Lov�����J���e�M,�{�in���}?*�/]=�T����������G�'_&�m������.Bg�,ъd�+�Rj.���}��M��.ּ����89�a��;ݩ�*N�ʝ+W[w�n�Y���� �M�h�tm� ��5A*6J��i�m�O���3R9kf��b?-��N��b�{E���N^l���U��>��*y�;�y:��j1��'zD�2̖�� S#�F+]�D���o�bw�֬��Y���K�F�ϙQZ��Ҫ�,�0╶K]��Ֆ��EK;��M)W�%�+��NG�i���Ҍj�����]�@�.�V)z�G��N����S6A��ז���B�@v��s����\�W���5t���|���Q܉�;u$�`��"۫�S��I`�+����愰]w��/�u�N$����]�C0�L������i�~�Etb����0�_��5đ�����6SS'ǩ[m;a���&�VO��]��(�啣5U�<�z��O�F �Z�;���5H����}��c&�(�7K�Dy�Q��A����|Y�?M�h�]��]�aT���.k@tQ7�Hս���!��hڙJ@��tMyj�~���� ���{^U�4`}F]M��Җ8q!a����]<h����.]�}]�q���G �ܑy��c��2���&Z����!�!;OB�M��rMR8��|@6/H1��&�ϐ��_���=x7f^�w�11������ܓ���8���ɯ�5���-�n\��R`"�a��6��X����xJ��A��J���J��e&G3�/ӆbё(q�Ͷ�_�8��i�S��Z�b�:Ӭ>�ޜ�B,_ﾶ�GIϗf�\W7��MV/]k�G}xh'����!�"U{�s�Gną!%�w�M�A"����B����\��#��Νl�R;��ouGSӦ�ŕ�İ*�GP�-���D#.�nD9N��}L�@�:����<|?���ӗ_�f��P���G~���K)�?צ�Jg����&��Y+�	�#b�7O�[��u��an/�
.H /�bx�U3�C���Ԑ�\�eC���ʉ ~mJyx���X��_��
(����s����p��l�蟇�s߇��c�C�KAx���-�x֓�#o��p(瘁Zr��>�B�F��r�������)�����0���<H��1� 7��� K0�Y?�iV�&�4�n��o`1�$îg���)����#5���?OX�xdd�&͗���w�Č���A�g욍��|I���ׄ��e7&�#���+~�$D�cު�W�C�]�5�۝ SZ���`�۱�"V����␙�F��(����ް��qbזW��vg��)*EFY�?!�:�Zq����\�V��1�|��B�E%���ڝOimq����?�w�]�UA�Zrm���@ċ���!�-��<���3ޡ�� w���'B]ggW���:�3��Q�Mz>1\9�GT*�P���+�S%}�d%R���^�N���8~
n���UO2�۲bo����;��C��{����O�YM斏�,�½�)H�b���\�X�mZv���q����o���M���t�ҚI����逘�炦w����&�\j}��`"ɍi�r1�>}B�� ��Sw{K�9>��sb�It��?J�Y�cvs���q�XJ�iS�:�^mЀ��>,����{�zH��Eo&�,Ɂ(y1������2|n�f`���1��������O�­v�,ب*�0�I5.�=	n0���8D1���)��.��V�\�ͱ�����U�B�N(����Ş�� �P�����}|�}�Aum܄��%j68��ً5�����1�v(�w��5�3A.P��'/\`��^A�s.e���A�V�zG������j�zt|�����H�]�c�F����ۥd�T�-�:��f�*Պ��ֱ>�yϕ_��ؓi��MQE٤I1by��'ZDk��y��i�%��k�0�C}�?�gA�{�����E9,�~v�<cV����ͭ�,��Iхvvw�"�c�����Xa���t�ڶ��7�[B�h�@�Ã��#�$����L�U��b�q������!���G�*�w�-���y���^���`�څ�����~2��u$���>�T	�ڧ{��>s�'|�b��
ǑMZ��d�R}�Ě�10z��y�>״������4z_��|![h�"�=��:�J����I����ڿ��6��X���Z��������]_�ɽ�g2�Vh�+ʑ�%���]P-���4�6��-8��Gd��s����M\�N��(koG���$���jCdM���V�ϡ\e�GG����_0��l.8�~����<�$H$4�V�N�b읬��&���ʹ,Ƕ)N�88/�������Z��ú7_����}���d?R���T��N�ԉ���b���'�>�w��ݔƒ� vV(߷90J����/�$l�(u������꧛����IO,��&�Ʉ�/�琿���\��(s�Q�RN�ء�y�����l8���o#���<���P�P��>Kު�N�lDy��ҵR?�h���n�
Bkpk��~��L���TT�{�ې�ג���{FT>���M�(�t-��#��sȪR�����x'.�.,*��|h�z����eܾq8K�+7�p?�h�`F��N*`��By����Den%Zh��,�
|�����V����Y=z����#*d�,/�����M2(�	�g�I"�M��C����%���wA4����d��#(�ѷ�m��/Ʋ���6��#�����Ru��Ø��e\/3�K%�����C��5v�a�{�f���qU�L�Q��LC�^����G1f�A�jʡ����qyLz9�`�:���oC���np�����[4��-�SmzPHW9���l�32s�.kԠ�2�n	�)W�u�cu��&s��k����1�l�P`ey܃"��ࣽ�wBM��`��Y6ʔ�7S�-�AhӘJP��r�5��G�\�	0�eAZ@β�>oo;��2JƔ p�]�I~���RQ$��'f׽�*7�\tT������i+W����%s�`� ﻍ�;Q:�]�]x��K���M��&W?5*T4o�N�4 ��\�Bp�z���] ��H�j�gMhg�B���W��M����,;x5�cU��okx���(giP�+*\qb)���P�49�qpn}꘹���
� ����)�(��xZe�%D��u���Fe�KF�ċ� �������O�%�BY���w����x��cP�Ń��A�Yim��h3H����|}7�Os杖�ݤc��ς��LylM�w���D�KE��h��b��/[8�t���<�`i�����Ci��jx���2�֯�Gy�^�J¸-�KB��U3����'��*�A=r�<j�s�Egכ*!�l�3h�6rZ�������3��K� ����Aש(&���:��y gT9�X���/
�	g�Wb�k�~-��y��=�7>��JYҤad�� D
!��',��f,Ɂ�Jm�rv\���a]O��;X�0����Ѻ�l�L��X�A���b���3US,<y[�=�������=gq����D���ej��Yo���Pҟ?�>O�"eD�MP������&�x!U�̂���S<���5���]�	��>`���KobP>����Ú��Q���RT���@���<��sSy/A�O�,��X�p?�a(��x\�9οv�W���sH}�i|���U��
�@Xx<�S�5��1oTo<m�A�Z�����T�X}�լ'ʝ���--��?��O&6�f����!�M>�"��Y�]/��j�q;�d�Zl�����[���[[���Q)�In����~7�%JJ��kr���yd��mȽV&���Th���}�������R��"������t+��t�r���ky)��F}#S��H�9�2�k�\�g.C'x��B9�ذ�L</٣(�q����>w'}	��;|d+A[�o1vdt�y�ߡ�i��a��By,�`AnfJ���;>5h�^�6���ŭ�7k�P�;���*���Pe.��8H��6I��xm�#��������CQ܀@6z(8�m�3i���s)��T%�W���ߦ,o;�&�9,�
��%���>?��
���$�@�y٬�r{Kß��i����U�����Շ�^��?/U 7�E�99�n���}��|	'�z�����dP|�PG�A�?їȊ�%�]h��tMv�{�<U����
T��g��U�)�C8��I�N�
 �6��e�s!��j#c�6h��h����C�C~*2f/+�D,�3����{p�ǃ�		�����������\39�?��ֽ���5lФ�p���ŧ�y�Mx����b�f-�=�[��v��PlH ����~�_�R�';k�R>'+��T�K�>'#l�6���!0�oBm�p�g?̕���Ĩ���Q�1�ʿߌ*�$�;���/8��Vb��~AN�RZ��6�DU����c���rS��i��rF���{ْev��Z�Cm�x�e�d�Jiy�- @־��c
߿�h�վ� t�g0�\ꩦ|�45�o^��1��l��I��qe@���ݛXN�j@E^"�v\��������ֿ ��7Q�[g���{Bi+_��R^�VҴX�B[h�!;(iZX��Y�Fz �+��JH���PNgK��*�F{�KI�.�oC�.�`)*�"�θb;�v���\��f-.����ޓ�ҡM��!���e��P�"neW�d� .��x�S���^�LB�ƛm`�L%{��rVf�.�s#e��y�]8��w������2��6�� ��{�$N;� ��?Շ��-�^��Y�py\�ɺƦo��d�]6���x\���(�ȟ6��^H�x:���Glk��������	�]?�&�*ja�D����p��RO�Z��v�&�u(�L%x��&��U
��ѣ��L2�|E��oweZ�����Q��i�i ��+�J
Wy�tH2���NW�er����V�ߟ����/x�V�g4j���˳c���;�`�	��}g���n���!cpʖ����+N"Y�q�p(R�nP������k���X���)��Π.���َ�̈��ܰ��NĚ~�4'�,P�(����03�����n^*=Q9����m����y�RXj�s����I����&*hO}�g �Gn̾ў�_��
��U'��c�Υؓ��Ը�eP�
��G�Oơ��^�ল1d��	@�ɻ���YY�e��jԊ)=�x�ڷ��xx�	^n9�恃U�'��w�	�F2�-�%܍x�=�I� ���Xl���V F[6�����b����yo������n;As��~�-��!�%y.QcV@�G3����Bӌ�񔦇>a)���y�9D;P@2F9�<C�#.2��q�c-N����w��h]��8�����`mNy��:��������Mى�g�I?�f���GS)��ON>��`1WN�('������d���ۂ�L�x��K�"���Z��3C]�g�:�GD��� KP8�ɻ�!�85���ʁ�\ t��e!ȥF����H}�}|侽H��*�`�����<æ�h���P�~�c��	��A������L�YY��g���*yk��^@���TV�l��%Iy+%�>�#��1w�_O([<��[��标P�\{��=3�,Y�#0MҔk�o�\��t�*�d�Fz,e7}3Zڥ��|g)pe�!�n�������垠2�U�sb��%��
���3�'�3d�/�pn�x�����"n:`kt��ʃD�Lpֵ�>�j�����Ã�&o�GS����݅��ӛ�7W�6�=m~�A�W�K矉.�51�-��yzB�-s��������"�������"#��4��ND�A'5�����O�uC:�� �X^�%١�����'TA���Pn����KOe��cN����{�6�#�bZZ���x�OvX��|�/���F�*����df1 �V��*�R�~���׹~���q�Q�{P���fȐ[���E�Y��$��ģ�̨���Q`�\����g�Q>/7���Ɛ�Y�2���
�@��$��kt'��S���	��6Zw�e]��bHBRD��~z��NHbe8�({�BPH}�^#����+s����yx^�l�U�L���^���%�+��b�a1� �����(���E�R�H�/�|�/��u�)���y=���_�t3/�'�Z~oCzȏ�O�|�i��#��7�H�F����.�&�_oOA(��vf�"�lַ(Qp��?�y��G��Q����%�oP"~%r���K�!=vÚ�����v}�@�y�޻|�����3TK9�dχ���F_�bT���b-0���=��I�zK٧�1V��u`�$J,d�q��Ժ[Yf���5,Yy��-���L�`C��^3�ڍ
<D�۠���,v������t�|�Ir�#��!�X����7�bF^R�@�����#G]ï�2��̯�lsQZ{�'a����7��M�G'�cR�:	��Sߪh�׎�*n:D�~�+֭�N��>��NL�ƀW�8�����bl���_�>�8R���=��v�s�i*z�P�I�0!��I�l^nU��%��/@�fFa��M-MWK�Q7 Ӱ�S��3L�'֨� ���f��kD��i�͆��1�b�D�Ƿ���bǔ�
�_v���DZ�?�G�|g����ݏ5h�OL^�l�?�Ht<��x�8�d�����>��/_k!�
GH��{�9�������Y�VP.�/[���3��Zu@�rƎ l�v|P�`S{I��b�8di��g��'m��j�.f��}Q���F7�~uD �V�`��4�x%�7r�:�)�#�C�F�����fW֧$Sp�,�!8�7�(BqK���^���^/Pכ{vI�p����x�X
|}^�K�7|Y�׫�A|W|�P�Y�t=�L���ʗ��<�fe�+찳�p _�/rlr%�{���������6Kl��ޣ��8�8i�c����I��c��g�3��|�]Hŉ���i�i#&�)x�Z��
aݸ�z��ґ�4�4�n���z3���K#+���=[xf�<�"n(Oqs�k��M��� ->�U�f�~;��y�%h }'_��p�T9�2���c��$����x�&޵0Ļ�g�FJ=��L�|�x%v�����	��_B�'3�����qd�ЫU��'�	��>#�)�̛4͎�%K^�Uff���6O�^Ȍbll��Vs��CUF�X�s�i0��1��W*Qf|ڟ��A`ˋ7WLa�����r��kq� ����\��͊"�3$DS�ޚ�7��+�$0��)Ox�g�Q�AJ�SG�=��{�U��������o�Y���}Ė'�֋\<E��6����n��-?n���5i_D�˒G���E�P�&��&M�/��Fs��{kS�ʖG	 ̾ߎh��G�ZR���-���/���ٮ�f�:� ��=$}E�$:7��T�i%fJ
�/t�'���	ZY�������po�+/��_�r���=�a3<�
1њD������g�v�7��>(�0!/�_���)�-�B5���:&D����#O��am�nE!Ȣv��w��O�]m��S����Yk�M�'t�E\�<H2�`ȕx?9�@!Ӭ9�PP��n���v�y8 ��_rVZ)�!��Wd)�?x�nOH�Xͫ=">]ʊ��\�s�Pv���p/.��j�3�(\���6w��]��/2�%����>	��d�8��R��5>�����6n�C�#%P����o�9Q���C�~~姧�u�]�sN�"�o0!^ł���ӁSfeߚ��a�3�sn�a�9g�2�[�VX*��Ar°�V ���*A��] �J�fOH��ߛR�2\
um��},���8ǎ$_�l�y�=)[�dN8!��<@��@t� Y�5)���x����q�޽�5K\M2ȧg*�H�&s�v��_s�����P��FX�#�[U�m:�@%!���HVOiDޭ�S��<�e������u�s����x�?/�PI�xl��� ��T3�=w���7Bm�v:�����K,�ryW �S��v& z��%fY��rU�i͌���&8Y��۶@Ia��!][�,�5����$��z��I���K�'�-�3l���:BCN�"�O�6=�m����ό#�����{�E~���L �ĜV�X��u�uK�Ce���� V�|���J�)�/����U�����m�x[�}�ok�=W>�L[*�����k��4�4������|M!vC"3���_GWW��Sރ�<P�q����-g.L~��*a�jB�}�Gc*�����_����0��:���2Y*i��u�~<=�^°��C_���Ղ�Z"΂
|�������˹@��>1��A�2ű�YI�[j�eJ����Y"�~��!��� Q��=x[������D��D�\Hݔ�6�#�R"��c�����R�瞧	_�l����J�� ���%;{M�ه�+FeQ��(�b��Eňu��V� �M��4�8P��:՝$r���c ������C��o��8_�X�(�Z�������LC���@����!�u�.t��Q�߄��F9Pb�)��{�|��Ui����v�V��&��3ٙyk皿�,�T�+P��f��h��尯`�
߳�/9��Y��T�QQi:t��t�R����J�D�FP@z���4���.$R�I���K )�%|�������9���^k����$���ah>%~�`z�81�Zky�mCb�S�A"�&��Q�}��X�s�B���c:da6�;'���	仁r&_�mtZ i��y�R��tz�oyNocNCE �����N�����qˮ�.Q�2K��f���wXL�$�/���(	����fs�ly����nN���f��~��wVw�3V�_T��$Fj(㽰�F�}m�/era�؉�e�iٝy.�ͽ�]ߜ�nU��Tjr*�;�poS{�ݑ�,�w��o��L��>���������}󻚝�E=~���ۣ Z�Ƴ�?�[�	� {Չ����P�v��w�l�e?�Z�B��/dKҺ�����q�3%G>�6Ȓ��-z�7��˔����������tlv��M���I<m[R��=����o�k��K�O����'L�z9+dO��o8H�.�3ջ�z��=9�� �읭�C)���d�5l�Md��UC��h`I���?�}��Pt���z��R�#�:'�1HU�[�����"�zI�xZ��K0�	�:�zݔ$]N���A�?��kj���=�K3DP�9kgae�'�<��#�t�}��6�@^�\ǵة\4�?Z����M�G40��mLU�koP�W�X�2���.m��ՅJ�o���U��	� �1"y��׋���?�j}�!�K�\^���BZ�4���� ��Y�>F�m<���u]��<ژ_G�����;x٫//
�uxt�4�M�7}����0�Y!@�yc�Vrd�~i������_��kpEs(̭r~~K��Y�sW_�����{���f^xBK�(�e�[r-��� VP�fbt��ѩO�]���
'
K���Ej�k��#}�>$f� ��F E\��lz���6��|�Ҋ���������l/U�\�NC{{��a�5ϛ<����n|%������$���"_�|UsW@���[�z��>��X©P���`��M��ȫ� :�#��'��o^�	�Ni���at]քpw �/!�L�z4}��oQ�O�C��e�5Wia����A��n�Pś7 �� 󰽠gD��b{�A+X�k̎�*���N
��C��=!��˦�b~�$������5���߆���9Z���ё m�ٌ�[X
�������gՏ�`��<�M	�:DA�-�N�7q.�� Ct�\[�����!�z��m*v�T<|N{��7=֓�ڔ�Jo*����!x����E��[��~F�d�t=RV(;�!���:���D7���j�<*	���Y؞A{d�8�R�~�pu����hQg$�iP�椞
		�X�G��
��L�b0y��-��fZ�]�c��7�e�e���ʓ���̲ԯ�K�z�)��R�%oٖٴ��#?�U,���o>���.�Q�W�K��������@Q�5�X-�\�ǲƵ40�]�R�s��,��4A��IC�� ���~G�������4Z�}���PM�:#p8�R���gb���F��?��oԤ-
���M�O���Z�X4��I�g:+��ku���V��(��[�M���Wy&��y��I��_��~��:&����R��n��u������j������Y�/�m��>=�6;��������+}�����i�u�^W�A�����4��Ѣ3玮(pe?Z'�u�-Ę�E�o�&&��BzA\Q./7�>�Q��%����΢���i@f{������7N4#Z�Sϐ�;��;���O�����DJ�?D�-X;���u��3�U���E=^N��P�j��'�g(ex��s��P�����@���L�/v>J���[D.�� <�X��I��b��̔%uH�S4A��-�@�;{���L�8��}'���I�����a&��()��+��.#N�࣏!�4�a�/H��d��j�L�+�JIg�*4t�0_dg���
��˂��9 �
5Mf�+E����=J}g�	��0��)�X��o��7�9Eu�eF5>t�������w��f�c�Iz�.躙�)��r����P�C���^0�����a~���x��pÉ���A���<A�[��'}`x����V�:y��n0/��5O�(�(Y���2�I`\�)���Oc�O���-�����⫱��,�!�~-v�h����3���h�_�|7 ���������7�`����}��л,��P��et>�IyK�11	3�rd��$�h3Lr�`�R���у�i��/�M	|{3�˳�������{S��9bO�Ob3���������&,o���Q;�Xqgv��A-/��~.�����F+5��l�k⽬����9/����Q
8�D������K�w����ţY�ާ~h�ʲ�(]�t�#�j�M3�Gދ΅sz���nM4�C�(\��;R��U�C��J�µ�tI�@1���hv�id��@��/�����ε�?_����Ӝ�n��#:5�g�^j��`V����eJw�� q��9,�M�r��}�yg�Tz�D3����w���N���e���۝����O���xa��Pe���<O���zD=[�e�S8t�`a��W(���j�q�z�4��B�f�L�&��J�֨�M"O���������J���A��[�o���K d@[���>T>|�f�%Y]?Kp�ZX+�-3 i�d`�\/i�\��*I�,�B��lG��	�{5�6k�WM����Q�'�(N�omW�X���_��Ԃ��5(Ri5�#��'V�?Ӵ\t�L.F�`Lۋ'zObRG��m�� �O��b�aԷ�������E�������s2!�"��Q4d�i�;"�^n�Ô�[i ��5=��p������dyI>kH,hKC�rڨR?�[����A��_�$J����L�&��P�Z2�Q,-������x�?TRx"��<�PTFwƽ�����?���,ZoC۲j��<�4���Eut�C�Z��?)IU�/�y�]����������8��[hlbR�%�j^v�� �W�c�:�^wnѥK�1|�N�{����THNb/>�E���n���p��i��W���؉��)�K�'W�[��v�GB8Ll����|��$]�2UP�����1Ǐ3*�3�wF\e7VZY�i�\���I� /�؉��@6���Qh����b���b��/C�ge���Uװmt����<��_P��+��b�{����0w/���oBL�w����
���f�U]��f輯�����BY�t��t��9[�� f�i���q�A,��w�УB~Ě��S��ƚ���޻ /��C�l�8輸� =� ��Ј�!D\J��*���TskQѤ�#
��X��t��Q܉����F,k3�T�W�0�D*��;� ��R���Q^���lʌ�@���_�!D	ǰ]��(ƲFF�B�u���;@�e�����*�s"�)c�'j�'R�2�f"v����Q=�Xg������'�����i16(�:���`��2
ڷf��Y���m��D	�ӎqNk����~:���r�����̪� ��>Ua/����d<�Rc���H4Bv��0�	�:�����؇��h�w�6=�>ZP�o���ਫ���,��sD����wg�S�`�U���_�W���$/��nx_^]g�s>��M]��@���bI\gQ'��,X�An��!)e	���x�.)���IN�ҙ�����5_�h:�
��5�g�M��J-���\u�t��*O���T�M�&~�K5�$r��} �T�A����@�j���Z����}��zNt�>����e�z#	���Z9e9�Y�]���N}��ÓL����u�	P��8���q>�?����nq����N��m�/��m��KK��0��C������1:�0�*`�8�JI��c��d�R���GZ�J�� �/������}����[�GY'@��������]�?�q?Ò^��T	�e���;��B6�\���2c�a��$�osA���x �Vs��`�3d#����)J��
5Q��_�S�bKt��s-���Y�,c-���'	?�Y)�z*���;~O��U��.�=�>��-�0�o�U_6e+(o����������j���J 1�[;�C�6J��I��;�b/U��M��fn�y�)h�8�)��GsU�b(�I�z���wO0���#��>��0��:�1�d
�QVo���<��J��0�?td���J1g�J��3~�^�Pzp[r,a��o�H��0��|�xM��Q���'+�d�Dae��w��Éw֙��S\��3�Bb���t���=	� �e�R:����[��0X��,����&��:�4��_>�ϴ1��+~���������-{���\�^}��%������a�;[q�Mާ��f��**�a�?EQ:V��@�gvg 	�'" ��~(#���yE/9?�t�t4��sW��I��(OP��,�Șڵ��9�c����h���X&Jd��7hꮻ���;�w���7-�{7�NU5��?�h�;ƃ�C�ט)�"�?\��.��o���+9"��x3�-p�e�P[+2w����Xǥ�EE�I�þ�Y��ׅ~j��3|m^C%/�������r}b{��鍛-�X�������@B�}��)U��j����
��~r�9;=s�L�Q
��}�P��p4�&��/6>y��
p����vX�"YD�Z�=�'P���WecT�.c�6g�zyE���\?ۺ�-jKVL��܋��W��:�w�H�?�w�u^"�xj�9e����+92O{t���sAa���+����gT�G)��~ "�t(��|~l�,���-D����W�v��M�Ã� ͋�u�e�k����	Ը�Gt���#m����[ya��6��K�!
AΜ�yNl5��R��E+-k���q�	��0��",F�o������3	$w���ZX?ؑ\�L.�v䎒��Q�;N��ʕ]�1[5kx.���~45�Z�-@8�r�/��o�u�A�����)\�e�٩.�d?�$��jO�!��v�;5
v�3��|�!����h�.KP@e�ak��Y0�3��y��dd/��=�|~�h"y����*�Y���5���ws���QY]TX��zC��m�[��V�tUO�8����fR�Dʹo9���O�	FH����`����[3�S�e�V���LQR�L �{����2i皩�cv�6C�'����{K�ۻ�u����U��l� ��U���,��{��XcO�~�!��!
!�D�H��խ�*P�Y{0�T+��K�zGO~����J�����n����K��&��o�bE@@/�
�a(�Ms JDw���%��z��M#��a�g��٫1C��+s�"{Zjy������O����
{C��${>�0�n��+]Yx��D���0�� C�Nkɦwd�Sr����:(DU�*����.O^���u�$ئ��Hs�A���&�b�_q��\��x9Y������?7����F��k�NlK�$`H�BRv��i���Iِ�t�~L|��o���Xߚ-�bj����r̱x.Q�R⚬�辡Ŧ)QH%�cY-�W�n��c%A��]�)d��p��_��9��#�{���1�uB��j^9�+?��g�wiP�M��	f�C]!9�'>�9+����[��S4I���VJ��˖̳T
옓�E��0[��G�Zԉ%N��yib�gG]�ǈ�-�Z��E'tT}�(�P��p�s^;���R�&*{���ÖV�y�����V�Iנr�FF��8��-d�:n��K�� ��^����>��ত-��9���7&16>y� ¯��P�5]x���ٵ �}�k����vRH��͜}�9P�/G��	�l�:<T=Φ���ߜ�h�������R�Q���3PR�E��kU�#��/��:���@6�c=�RO�q76�K�$_�U�"�U���L:(�6,�'	��s�[K)���JOJ�a4('K�E�b��2������
�£� ���lcR߉w�HH:�T�^�4�)�|}T{\��>\�ys�l��5�qF�SpW�%�f�['Q'3����$ϲ����'ӷQkQ\�6< xْɁRw*�A8���\;p�zy�D 053)�e��2����h
Y����B�G�?���Pa)��zP�Č�_t��N��ݚ�PlJ��*��p^�P���c�'� .����Ue�3�Q�k��2�I��V�5ڥ^v6w�z�r��;��v©������Gɑ>_��������M�)�j�o�����ܚ+���O)|��}����5I��(�xb)�@B ��L�p��,��r��.V^��0���+�am�݉x*������{n�F�߲��)E�\B���Ⱥ�>=��+ɛ�I�t F!���,�����8^a����̖�iϠ+\Ps�I�l���%6zA�45�N��2��#������-5J@SuH'�Y��B�vy�Z�+!
��@���oe�[�e���)�����h[�D�Џ��,���)�'�	{�'4g��]�1�i�ΙSAE��	~�x����DV����U���`�PjU�y���P?�� <��5о�9��?�؝��95��Ѳ#K9��-�&�����\�y�β�=~>��~��4�7�(-ǩ�q�9�f��[��^�e=����b�,<�����1Q�U�3�����̓i��(52��/f�_k��?cf&��y�Ƨu@��I��l0��oJ �������i�Xf�E֡+��V^�ᤗ+*���)m�@Ŗqmƪ����v�7ր$�B�S�}\l�RА
�ͽ�~8h��w�v�bo�m�w��n=���
�{���?�7�j��qG&Z��s-�S_�1���ǽ_��Dz�E�EA�V7+<H[��9v�l��
�f ըV��i�s:_�e���N�<��w�X�ǽ��j���A�֜.t���OposS*ң�y~��;���e��sV�6�țՆ�=�O�	�fB��l�d�����{K��C����� ���gƺ3���2]cV��Y�N8�D���>���W�n����)[��2�.A]��#)v�����
��/��=0lE�3})Hi�GDPLh/@�|�x�.���I��IFgA�X�����`�SE�=�U�Fy�qؙF�u;��}��}�L����P��PV�H�)�}=J���_���*��4Kɋ�B��^�+{Y^R/��[E��Z��Fl������d�,�'�w����2���ki��,P��w��6*$��#�i$*q)"���z�?[X���&�S2�%~�{غ��KI61�n�6wV��������.�����V[7ބ�f��E�	@�қ��!��Lg�?!uPG���di�q��o�AS@;3�Hac/g:$z��r�ϻ�����$~X������(�n���V�gp�H�(��3�
j��
��AG��ӄ}�XpEG�L�E���=��&��T<�iX�!��	EA����.d-l�^e�z6H�.
�[���o��U��2�/���@���F�n�>����4��K��8f�2�s�=�VY����i�KA�C ��ӥ��7��Q3aSR�c���
0&O4V�q�� D߄ڜ�����*��������ד ���Е�:5�����2��j�BP��KΣ����;[oR���'�uzԦ�͚��(u2fG���q	�EX<��{Z��� �j�e�G�.% ��Iv����;ң"XH����h[�e֝1�tk�S�p�::�ߪ?�X[�)od��_߅&Ph����6�m�#�[!����Xhp]n��^�%V���Gx�ᶽ�_-���.p%6�ڢ����p���i�S�V���[:�	\s駷X=�)�J?jQ�5�� ��\��1��
��#\�b��qɠ��Y���d0-���X�߂~�5a����̭��M��1���NvQ��ٿ~�9 �ײ�;,�%�i-��
j�u�bs2��ٶ�v�O���d��O(���?��kl{3U5�p5�]0����T��|Cgr�=��{�JƦ��{:r��˪��ݹ�i�)h�}́x��EY��0���zǎ�L��%Yc���_[]��p��%<��0%:�+��V]��/}�!�G5Z��i��N�x�`�9�#w��Y�d�	�'6���7p,����;���jɴ�T�v�y5	��̪�	�qăE���h �����]��� i����=_Y��"��T>�%?�v�Wm3��c�fb 񯓎�����������0�d`m�f��k�������H$'��Gc�g�u��Y��iOj��ɻ�#}Z4�%�>o��M�R��71õ#�A����-@d����	���-���&��t:'����2�[�I?��grd��o=��H���Z��ђ���h��K����E�0�7�$+�4��E�-V ���~:.W�2x���	u�������u�%4�
���)M�ΥQ�'lv�)s��ƻ%d�l�hsL��=&:m=��������}�&�->bxL�bטC�jNH�kvώ���+�_+)����c�QZ�=N� 9�!�8M������������v�#\�%+o�����8k�ԩIq�R��A��A<1�=�9�b�*k&����G^�N����������fV:��{L����@F������'z��­p`J���9_�N�]w}m��|��7[~Wa��W5��2&��GU��|�/{q�Y3_* �g�`��'��>Q��nVv[���t(O�%:�i:1�S�߮��N�	�����8�
��X򧝯1$��\�5��lk�����}���_���q@�ݦ���A�oQ����� �2=��S`v0]��;�3L0��6�x �A�R�Y`�d��3>�A�|��7��3��%��1h��:��kwxBk�ѿ��Z��+x�3������lp�Nd���24#�x�]�Ɇ�6Y��D�T�pl�E�{��d�Z'b���������;z��T\��ʻ�'��?� 0a^�eA���Uh�O��4�3����`k��{�9�Ԗ�q_jF�� �2'�
�%�'�Td��jE�|F駟wm8��7��~R���ʞ�㑺r���Ɔ-�����~���|���M�-M'Kk�M�0��ޘ���z�WN���HW�瓝�K}gn��<�k���~�.������u��O�����XoZ�'�^@cG�J4A��!���-��j��N��A?oɣ�ki(�32��9_�y��O"M$�*	����񯙓&�Y}���qKͫ��2����pz��+%,7�����$hv�׹���e�A�%�;�*���!D�z�y�
LX������k���l>/.7苅���=MQ5���E�U���_����+��^tԜ�L�G��K��uy:7�?(ނuE�D)��5f�v�ǉ}��J���t���5�ܑp���[�vhe���M5wr�Xo�O�����'�9���'J��d���Z�j���ߑ_��s����̍wP�)p�V��.E`����'o�'d�����Չ��O��+M�_��v�	z�Aw!�g�ȋC&4�v�Ž���U�tq�sЗa�� MM������ms��<5M�c^O��=�ePg�ԝM�֟�3�T%���ى>�gA;r����_��oX��}Ŧ$��γK��xC	;B�h��9(�������}�/a,	g�)��(�(BW=w��ظA�D'9�ĜOwN�۪?Z���tG���L�h���갲��C7��[���Z���+*�%ɳ��+{U?�UW5�M5Oa�/�`//*�X�+z#��!8K�έ�1�j.{%.ٖ�x��܃l��F��z���#H��Q�~�56��.L����jD����l�Bu[�<�~��
���!D�T��\�g�tl͏�>^^2��2��Cᅁ�Y�r��@�Upߵ5�ݏM�l���(���c|ݧP}�
ԶG�@�X��M���W�waH�Eɷ��Ϊ�x��"]�N�~�i��	J�|�@.��N�"�=�mM0�nk^�����^�^<\ �a��O�_�Y"�����?� @q��ٽ��Y��**�9��b&��z*��nL�t`�@�{8�沝�?/����?��8�I�J<�1�A�\��
�J��6�k5�`*�t#��6���|n}}��I�5�����|�7����>��$��&(Qu�a��uh+h��=I�Ϙޠ�!�|
�oR.�B-�Q�C:-�C5 �r��WJ��=�d�*(����u%�Έ[7�շ�r�7P�0G���f\j��q��+�����keI���=u$]t@�h��
�X��b�����ݘ�ɝ>��g2���k����|3H�ZrE��1��c��߆WK����h���H���c"䌧�q!�)η��t�'��P^l�Z���R.ն�>O�F:��??����AKy�M�6��B��^��?-��n�$*:��L ؐ�yd����vA��#��,��i�D��f)�{Sv �k^a{�T6��V!�VGp��b���]\Й,?'p���=l��w{[�.c�Z��1��^K��"�tt/tQYWʍΦ�I��M�p�/H���!&�m�lg�'�"	����+� �:���F\���c[n����n[>�Q�\:u�5c�
��M~�N_h����|�?�F���an�\���N��ә�@P2?R�m�tx
&ٿ<��Bk)4�IOs��r@����:Jr!���Sk����$����������v�h����l�r�n�I�u�S��V��).��L��^��y�y���먨�*�Ç��$��~?Q�6�L�o+��A��H&�5�t����k�`'�u\D:h�u�l �z�� %J4J�u�����-pI��j֮��Ti��[���p�2�4�~D~�&b���Q �^?�:|�4:^����pL��Vq�ej�� !���03���z�������A#]��^'�\�.J ����|0�ͤJ�p����'{|`�7�H^=�4&�?.�p=�P��m{��t�-u���$�/{�{��j	�O��6�+b&L�S��Z�92�,2��Y-�b ��p'�����}FX�9��'?��qF�(�c_)�`�:y�#�^�A�8^�;y��
T�F�UX�]�@ �n��cVҗP��)u��4��:B���0y7��H��~�l{��U'ׁ��!�p(�{��UNI�i�ڟ���T��y2M�#�(D^���/�z��柘9�&b���Cמ���jo�$&��mN����)�Z˃J��������Zd����]"�A�q���fW��:s1	lÒhe��	�[�i�ʖn� b��:��F���XxV�F�*��3��g]^��rX�l�MdQ�����voU��w\�����Bo]��sVU6t����� �)/R
㩨@�0�dd �Y��e�f"�4���{Y0�h(f����m�]��ԥ�Bm��B�V��$�G�#��&��9���2�0ݸ�Ǣ�f ��׹�W��ֿ���G�L�%�]��d��G���7�����T :*�b�q}�.tfV�R�%鑝;%q �vzKw�۰=r�W��@�d1�U�n�!�V8\�K��P�S�����y�z�#{\�0���8پ!��]�&r�ӓ�0�1����B��
s���E�#�\�LU�dʲ��vܱf�:-uHBA�O��Ti�5��`�G1����}R�.\2�Sn��j�Bz�U�m9��_���A�n��B�#���p���������*y���"2��8�AF�Ic����_=;}�{fe����*'k���$odU!,!96���~x�o�T�����J؏-���~1��q:��5lվW"5���I�������%˝�5֕&���]|)��%�c�-%ک��I�X�纶��$�:�f�t��($:�v-
�N�d3�^�9h݋3�W+\�ؽ9��<��s���7^3,�]�ai*S'#1�	�����;�.�h���c(&��c��� ���ّ�Ed�!q�o#9g^�}��>p4HI�0�C�l�gK]����������o�Ő8c��S�l�In�=�[�gh��k�(�iV ���?8��@�Κ��{vƏ�o�.�|�����	��	Ҫ:�����j�2��x�[Ԣl�����j1[���W�����X��k8��mޥ�^:��EhQ��/D45`.�$+���d�L{�a��|va���yU��`=��x��$����2�z� � �	�Y��%�#��6�ug�j�ͦ$���`�b���g�3f��\qQU��V7�Y{>�5�oHU�]� o��e�h�����5�h�z҇���s��_��9<�c��9� ��H��[Ma*%�Sccr�GH�^EԿ���=��s��>���M�w�� �Ap�j���'�����ޫ�ݸ4�,�	�N�T(����%���c��k��t ���M�U˷:���49˖�ǡd5��@��)�J;���?�J ݗ��'y��B��u��]��r���-���p fQ�UȦ���A+�Z�jXi�I;� 8�]Tn�Wt�J1�1���b��^�g�D�7��[,�S����!59��$���"��}ش�Ŷe0���\n"�H�|���XzS}�^���$ɝ''?�II������8��R��,S������(kÝ�
+|�Vk�Z��!Q��T���,R���V@>1�ΐ~��[.t�Zx/�/Á���������D`�w�3���n_�w��x�p".�Ua���׃�lY�Å�n��-�����x�x�d"w4~Z������iT�˃o�uS@gu�#1N�{�ȁ��Cꄳ�C,NP̘�Cαrs
�D��j���4��j%��χA/Ӏ�-�@��Y��UB#�[�XG��f�����.A�yA	��웱����by�Dv�Ļ�*_���LsSs�WA�(��'�><����kY�pS�Ę�
>/��Gi�֢=���-�Ŝp �ZK�.#���LS��J�+Ie��g����� �a���5oyS»q�� rd��<	z��k��ˋ�}WҶ2&~@�W T��re�qG���%m�=��\�-9sd���.P� Օ����ݖ��˩���m��(`�A�7#���(���Ts�+����Ӡ����i'��%��_��\c�	�u��z?|pMb �{��|dgQ1��n�S�U�6�y�͡�KY���v�N>G"���W�^�0;!��[K^�]KlT*�$Q�z�O�Fl�5<)\1P�s(.�w���[8�Z���t�e���R���Ԯ�`w'#�,q����g��t��V?�4-�f��kr��NOP	��Vk�NP���(S"��pP�t%)L��Ȋ�&��d�'��}��7g+�Z�r���6��.B<t�ZS�\8k�9C�#�`G;���e��S��*�̇ug�d���TS�h�BL�Y0�'�3����KE�P7=XJe/��O��)���c���`����J��83�j�>��[9�M���]}�����﷒Fu�n�oap�Qԗ5A;��ih�Bm��{K��sU��<_�������X��V1
���Oj�7h�����plݛ:����Gm�n3'�ř�;�������k�j���y�g�`~d�*e����2UU��X�ޥ���(6��Nl�Ru�����c�鰙����,3�ga#��+�;��y�z���,0#�;O���ظe�L�Pp��[�v천ZX��lZ1`�@����;�!z��6\�6/J�c�@}+D隷�S3\�ރ�*��m�5��:J7�a��f�*��Y��۱�O\�:��绂�F��v��Ƶ�з��=`�#��|j��}i�l�ٰ��������r�����o �%|�� aw���f�&��ޠ�6�hԧ³<Et3{�䩅cej]tw�}��ݗ6�߁�O���	l����G�H��) �yx�:ha6�q���p�/Џx�ti����%�+C�㯝�RҰL��<��ԑݣ����3Ml:���*���ö(^��.(������_A���)x�����j��F��;����s��?���zg��R�0��d/δ�K��ޏ�� ��$�`i���=@}4��wBӔ��;�3]��uڥ�{a��>���(��`źϘ~��44��`�l L��-�$ @4�G^m0�	�?{pf�eZo��W0��:Tc�)3��RI�V�t���ã���.�:O��$P(��l��p%&{P	�$�X�h��O�h�����:,}=��\($Sf����4���ͱg�Mu���Y�Z�
�B\_���a�R�T�����C�>[���;S�.Â{M�����@ն�D`�#@!6&���^�ٟq��E��L|g��u�������G�m�#w긁����t~7>*��"�!�C�J�٠5�h�e"�d���u��nZ�P[���(Q��7�e�R"Oq9y��h)=.3��X�j���VaVCO,a��@�U��1����FW�~�fml����, y���\"����*/s�`@��?�����~���Ğ��E�l��5��i��y_�Z�[�[�Q{��i�`p�%�,��k��O�'�b�?�����m*�3���4�P��px�-cB�`�C%Y7��P.�6d���ii�d��Xa�j"f{.�2*�\�l!zl�@p�шPdȐ~��2U����d����+�r+\��J�7�'R�ɬ7# �ԅ���B� 3x�arwTF?�_u���3�5,��]���0��(_�V���l5&d�G>l"�#��~T�q���x���^5�x�n���m���Ym����rhu�r��h+�6�.��u���~ؿG%`=l���ƃ$VpE`X�r�6ݠ*N1K�h|�YV"[�U1���� ~5�~��G�T���;�;�o��Ȑi!$�Br�n��ka"�x,�u
��o�V����㋼A�!�bh�9�K���,����F-Dsv���@�?�a9�`a�[n�A�A+��������[�.K���$y`���T�RFD�8�a��:��瓅���'�ٰik\�y�ߴ���B���N�]�ĺӃ_�T��	��np���*^~�]�^hL���z�K��P�5��E_��8�!J#]�#%��Ŀ�Y
Ԕ�&A'�z~%��$���9�I5���zHt��Ϙ�b���)��%�G
]x���/|���Dfe�m�c��0x�jbx��<!��D�p�+z8h�$2��Cbh��@H� ɟ�޷�íd3"Τ�'��*z�:v�e��:����]��^�z��Bvu���(C��pF�*��d��*(s4��?;�	̅����Td����iNM��K��9��жTn	L��mY��
�L����)n�2��]y�T�׮S��(�h���#�m���[t0Iş�\��3XG<S���rRxI�^���.A��v�Md��]f�|�z%�3F��k(z�����q�D�-�nS�_e�]���D#�����-��o�{;����7,0����E���# ����!J�Wy�����
��'Bx�E�H>JC�d}�U݋��B\xۊ�SAPJ��FD�I�/�`r�5�.t�<��o��{�f���6	_빺H&�t�di,�L�V,���$�R���J�#r�P��Ece�6����LdW(:Ȁ<sj�:H�-�E�����������G��}'ipJ�WĻAS�k3Љ;��>�/���i9�;����~�_�e�7��T����e���Ag�Zz��C;�����U���Ȕ��|u�me|�r,���ɼ+��b�R���>��@PP䫣TM�X�>%� )p�&��[$�����bH��|���L� ���0��@940���t�e#���0���W�޴;�b�)n@C-�F�Zg�i����I��W� �ݘ�~�&��)1Zn0[D��L`��|�H��נD�� ��t�!W�l����*W%/ J+�~�������(�{j��z��}Q	p��ow �Z� '�33�`���FYafZb�[�)�5�ٺh��SB��"^�9%R��T��j�j'R:��l�D�c��(Q���������!4:�g����Z�� �2�\����:9�&��MGJ�&�j#��T��w%>�KW0�.��6|�h���?�O�P�&���֭]��~
���m���jP2Y�g �y�mn.��d=�`�]}
�S���5�_�#�ZX��΂U�֟cM�K���3u�'��{���֌fb��SnZ���[�=V ����d=,M���Æ1��pGȐ�)�x�e�4�њ��{�W�w�\�ϳ%��5���w7E���,2r*ѪE�m��l�d��rc�Ѱ��?��:n�I�z�����Lf��Y�ގ(�\�W�9��gU
��J&<�׮F�S�#Ug0�6�\3��YN�/�~u �"�d�`��SC�s�;����.�̺Ш��U��xS�h�\�H|^��^��޲�q��EYU�G����iN0Z�9��d����;
n���!��-�����Y;���ZN�b�˞������~F��+kpWB�m�o�`�� Q&m}�x����6�ݖ�h�^O�������}%�(�@�j��V�"t#ҟ(��f���0�(�r�dQ3�'��@䕧��U������|�y �-DΣ�te�E"'��K�%�/�af����z�ϛ~#$�!T9_�`�P8�i��r����)�XZ�8�8~H}�DR+l�yj�t=��˘�t�eg(]P����B��-��\��G���+̪���y��yǯգ�-lG	��Ô��U 	�B'��a��Ma1���'��'+LM~�3a�Kqw����%�3�����Ǒ
��ҧh`6'�`6��:?`
�Q%�������xXn
�� �����C
�&���n���JR̈́>dc��7��-eo-͏�n���5[���c�s�2��E�'C��ȏ��{2��EF�
�O٢��ږ���h�y��w�c�_��v���̢�5))��U�ɺ�6$����XM|�m_�L�/9�%�>�ɼeN�cr���w	o*úL�!d?��>�қ�z8���� t����W�@cQ�z��\_i�q�wj�.�[���t��8�>�BpdXsX���B�OV������sv�D>j��M)2*%#�:�Jb<��%@���ٲ�v��Ւ�v�у���/7���98����ߺ)XL�^;����� s�:ȧ���	�/!6-V�@�\v�z�ޕ��͂k��o˨� ��jD*b���vߙ6����P$�w�Q�A��ڻ��:KE,����hn�)YF+Y�]����ɴLG�6�N�չ���qth]Om�E�=������R��s9��1?b�)f�T�c��vy|�W3v�a7g���K�W��$�[�>ls��@�FCLE�#dlP�&_��27Z c��YH��8O������W���W;����f�v=���X��D����b|����u;Ѻi~�Z��R�n�ќ��V*,��g�꠲7)�3t6�����	��k�o�_-��~tR�h<�v�A�����'�	>�ڵ�}�g¥��~�~��X�<���ڙ�\�?.�r@a)Spٺ��#���\��񑢓��"B�NI����rt({ٳGQ����RYRɒE�=�n��,��>�샱o��{F������龯�u�^����|]�}߳��E�jVb@���'��=��q;���$=# ���̉�vLk��evy�h*`0�O8�g����6I�S�|���q�ļVK�6I�0���i��^a�ޭ����?NRʱ���	�����
��4.�0�7�&�k�:ה�T���z��қPC��tJ������x>��>�-���G��l�?����M#���.��"V����v+�۳���� O�+�x������1��ex��j��4a�Fe�������)G!�Ѷf	���:�v����!G�w̶p.S�K?M� �Q���"��@�_/��`�c"�\���ETje5�fs����?���KA�L��P�Dټ���/��q�t�餧�}~���E���~ �
Ц�� D��f�o�MI�/z<W�������Z�I��̲f�y�eT���lwΖ'eF��!�>�T���6w�N7����_�u����^�q+'�|�����`"\��:�9�������0KO����n�E���y7��u��v��S?iju�z��KL�^�y�z�v�Qc����l|cOu)��0�'��92:|����ޗ��S.QW�ٌ��L�.JT�Ga�/�[�A៩~�v�ZP�1宫>�[�3�,�H����ּǵ��1t���`Ƴ���
i��� ��c�Hy��{�� &�O46j@#�{!���9=̧<
�2}��9�>Lw�=j�R�Ҥ ��a�2�M]�G5�\>g&n�`��(p��.PO�o{9宽�c�Շ'A|��/���/#��E�f�$���β�?}.��n���l��)��GYK�-�G�dzKΣX���#R^��?4��j^a���u�b�ř���J�v�O>-���_�̒���j�L��S6��+r�:X"�!�5旑���Gj��wG.�t3\�����{5R���ܞK_�-B�&;Vg+�a�3U���hk�r�e�2�Y29aP���z�3���N�*�4��Ԟr� Z�$�q��c������%�6�s[��ɭ.�s�4�o�o�;�~�ϳuD.��Q(`K���+����.�%�Tunvx�T�'4�A�d�c��<��H���S�-{���j���e��<������^�}t?#c��n(�?m�G�QG��^��Cv~r;��Y�����N�E���I)�3��r�<υzS����A�_ab~����W�5h�t)�7�����~��2;�����%rȖiF")#֡��'�+[��Ҡm��j�ԙ6F����\z�_�F޲��-*��!EUBB�\��,e�^�wi7�ps1�O}���B�+4�?�a���Cآ�Y�X�_�2w �Q�3�Щqk�B����Ϛ���\y��&e�=�C>�m!���+�a櫕�zC����6�c��9>��`��u,ci0��ު�Sm�c���O�JwNk�	?``�7^Έ�\�;:��H*�k��ut�H!7�F7�ӕ��7�QS��V`�R��^�:��,���cH�g;��_�L޲M���;����`�y�f�߯m |��j�8� ���������c��Ģ�a�)<�'�N������ ��w�Gn�D���O?��U�Ö36��DM��B;b�,����=�m��td6�R-Â�3]ꮏ]Γ�y�W0��I�P�V�'��S�A �O(t�5�m�+w_��*�,��[1%�M��Ѝ�_Ɍ�@�8��c�(XϕGH�A�����8���@qN�w�c�i���%D�PU����
HJE_n%o�-����+��w�@�) [@GD�%�N��u.��R���.��µ��E��s1���Y�K��MN��`���3[N�W�(�S���w�H^wד݊��]j?��J�ln��K��(�Q�jU��m�ݕ�1���h���������X�09�ݗ�d�C(�=���[&%3lw0��l�"�����ur���7l����߹�c��|���(>��S�T�#ڮ�n�n[���n1�CrG�*f�j�8�.8���5���b}�8o�/���%��_݈R�6�L&��2ϼ'�R�2,�Xr��f�l�cҎ�S�%J5w/��Y�2;�[e�q���5-~H[T�㿟@�csP'�|����:|�͝�]x�A�k��CfԂ�3�W+Z�
��/��ܓp�M����om�=C)��(t�AD��O�<�U)#���lE6�p���/0��(X,��Ŗ���7��kn�q�z�� �`;E�+���;�������*�5mvc�
�!��&D�cu�r�/�SID��ݼ�Q�߷�׹>��U��F��'��?���$�z����[_����m��s~#�5ɋ�e3,�%��5��q�A���k5`p�� C/uq-S�oѨ�_G�e̯_�7�F�Z�/E�Ǣ:�~B`E�}R�I0�5�E��?�ڑ��Zj�wɻn�Av	��a��g���y��Su�f�^Bgz[@�Q�����2:I���i�k,�|0	/����1�8�����4��M�}�r�Y+�U�C����(�� �^5�������7�P��x6f|@�n�L��j�F��龃q�����+�-=J$�ti�:��Gh��k�$>'i�D��.�n�����ޖ���R(=��˭:��Y��6���Ȗb�!8ws�����#��`����Ʌ��͗7l*�gq^i���X]�b;�ǵ���2 N����+�3b��J:/�Y�8�`��0ܥj��hG}�(�ϋ��r��4�
D�� @Y�	�zˑM�ۉg�`����܄��ϴ��Νp�\e)

A(���Rs��xy�w�V}��x�6+de��LA�E]��b�V�<�׏��X$��fͫ�u�t=k�jϽa���7 �mnb���ڒ���wz�S$x���>giH���A�.�V\"t~C�\���e����'��%�2]q������SW*:��S6��U�5���-|H��or��_�.H�����
��E5Ϭ�����F��n.·^'d����zK��*��3��u�<�soAM˿=�g�: (�7��ߗ�/¹�X�-w�
#,A|#OEM����|�x�+�V�d��T�%���F����?Mi�Y��;�_��G�T����QVS+ܝRX$l�&���
�A��ԴV36�*x��G�_���_���TP7hud7����z橥��Xt�����Ոpa��-t�J4'k�26fo���V
��Tq�P| ��ss!|���`�+@��o:P��1W��9�� u�Ÿ��M+���-�}D��V"+@�	ـ��9`���o]2����߂�o��~6��K�X#�֬xJ��Aua�_�p��A<�Q(�@6���B�(��^�����Ÿ�e>c�>w0���?����K�Z��ѻ�v�K���<0��I%o�Yʮ:�$�vS?�L͍��0����ާ�7���$���t���t���S��Dg��գa��T�z��=]��K�����<,�ɬ<��ۏk'}�1�\n�J3���9�B��f������?<���Y�&h���H�Ǜ�b���Kݑ��֭�"�����١�.�����ذ��p�qWש���w̫�ӿ��7�����}t�RJ9�E�C�M�C�>^@����-`�)og9�`����W���g�@�n�pd�ޕXɱu��=�;��3�/s�ҹ4��Kqgh�����q0.��C�DK��~|K����G�7�_��8e1�Ov1���D�ׇ#�h�m��Z�5��GNF-dAo%�7��e��Dd�?�L�6����j0��ODy.��Z���
'�ۨ��1� Y��x�^P@�f��a�c�5n�H�_�$�m� ��,�Z���K=��Y�d�zc(I�k0N�������C��
c����B˩��W�˭�'�#����(�mV���T@��#���o�p;SQnc1���*v���W]�]���/s�����\Y�l�����������F��ㇳ� A���<M~�N�^�a�D�g�1S)t��e	�zJc�'��
W)[6ײ+=E�F�'D��vE+	������=M��������j���UR��;W�=�)�2�k4*�e�4ʂ��^D�VEF�f�?���1��9=\���h�ظ2j�Y]���J�\A��2.%��LL�\s(Y���}*ea���L-��=�_	�|�U�y�`x?Hu�./q��+���Z'+�I6Jo���!XB����i�Ն�����k�>M X�٣��4C��s� *>@��PWX��v3��Q2B*i����CD�bQ�� �p��RAi��(?2�x���K��U��#��4�m��ʁ�t��2����>	C^,�hh�b;'s�(@���������D9٠�N��.��z��=U���qVWB����h��҃b>����e����s�K/����洗��o=�v:��$v��wr&z�SJi6��\=��}�'�C��q������)|�����,���ۏGI�˻�}
���&��G�I#��,�����Dߖ��E#�o�#�#]1��y�2V��i�J�13xS.�A��g�Ұ��M��,�:���Ʉ�M�	���ȃ4�|؇AR�,O?�u�hkQ{� q�L����-�q�,׽�=/�jH �72��s1ȇ��dbV����f��T���ҹ�ֺW�@�e�4�;{޸t:�]s}634��p�ȫ����})��3 �"A�ܟ+_,�ה�>y�B�b���{��u��bj����~���&�(P�_����?�ʻL��8��kO���xZ���z����X����4�	>���​�&�1��NV�g�����2ͬv]��0r �&�%f���}`AR�,�r֧��>6��=,yW)U�fn�^$�*�zو��wB}|=�sAw�Y൏�8��Ct��8����ՠ�v�����\�w��﹗�>��l��#�_�����R%��1T�9���9y\���/���4�uKq�@����[�k�����Fs��}���|��JA��bV*5ũ(�5��;-��!;a��i�-~?���'B�1�\!o�s�69<�w���4�Z~׷��pާ�X�+�kx._wA�"Xk��I����5)~g@N<�+��kh=��1��)�e_j�2�y��K��A-����s�`�ݹ����	� @{� �� �{��$&��� ���5��:QLn5�G>�1Wo�yc�?E�c���p�hF��*\�����K�0r����R�y��v���R*���gy`����ē:��9�oB�#}�M&�щ;W&Ke��vJ0�.��6���P�7`�o�V���ɬ���R���2���~A{���T��"�>�J$&�ށl�g��@4)$&j��_"��h�!�A�kC}l��M@V����*�c*�U����*ZL�~*v��ZII8�`(k�����ޡ͑��AsP]������h���p���պQ.���-�Wqi�,�q]CWҒ OQ�^"_"�Dx�kw��,u�zD=���`����qX&�9����8�y���a�B��qB�:���U|��t���E��70@�e�(�9�S�a� �fG2U�l#��7>�9�����sEf�R˦�,�z�`��}� ��#�|��Ј�b��� �>eu9*��]Pv�wr��s����za��Z�z��P�WcYŌ���8�<p0c��N+:�LN�+v���g��g���Tmi�0^d�{3�Y��a�SL���I+�	�6,�]#��fI�'�o��d\��b8@/'GTV�&�6�'��0?!R8���Sf6��ٶ
�y�����[_��L���I=��Ȧ�B�'���(:Z�E~} �t�Y O�h֦z"C���̩_�����C/���X�+��!TCq�\640��z	�Qm���	+w�2\�޾}Sv�}4+�'�9O&R+7�W��7!P�+�r�'E��m�]%�ͻ 	I�k�v�\
.��B�F���	��E����aH���_\
�;�z��@,�������<n60]��~���p3'�/M2B&�_�=Ȟۨ-c��i40����w���=�FI�:���R)�\��{ݧn&�d�`�T�2|�}�O�>�*��߱�c-�O_������M� �:Y�����ά�8���tI�/���H�*��ĿM*eڞ�^E�_����cjFo��B����*��߾/Q�DJ� (�˺�l���^)�Lt�v�~�>��:E\��ƀ6z���x���b���`��T:��n	��U��2��A/�k!�5p�	\���m|������5jI�����B֕�]�ݟ5��$С@т��H�P���.e� H?d#��>�m{��}�K���ry��8�D�嫍OT�aG�$ř�+	��/�rB����gxh�6X�|�j���db�ξ��II��C�&Þh�� V�4-�j7V���7�����ů CB[;�F�%�Ȃ0ˊN�<���}�Ӵ�e}U�ؗ�6A�60[���}'�&��2��nN'A����#�e'�e����F���=�m��h���n���{�F�Zo����h�=��!�"�,��=�[��֤^޴)h�����E�1���3�k�*��[�m9T���}�g��ۀ޶h�w��7P���:/[���2���ֵ��X!��(��*��!�	BP���2޴~M�vxM�p#�8��W��^ؖ�����[����S�"т�qz$���j��O�?�-��3��̣�m�L�t��
],Xr�D�#*S�Tt ��!Y��lu�� f�~�²�Ke��+�>�,��"���Iqz�Ç��Y"�ȶԋ�=��j ���ҿ�������n�}�~Kp����߫l��M�+Y����d�kD�r�J�K�j�B.�HɯH9hD� ��7�����ؕ7�!QG����X3�h�Ek����so�/�8?�@�j�5�.�=�a�~.��2'ʹ�VIKM+�;�XX`��9Fj_�(�[�K�L7�(A�c���]��������q���Y�fr<��9" >���f[c9�������W��z(���)P^ +e���\����
0�F�ѵ�&~��0h8(?p�"Q���	ӸK>��2kv[�er�P]9P�E���bt�\n������8�L�9����˼G�4��� ��̓�^��w�Ӂ_���bS{���/�!T��Q@�({H_�m*0�}&�d�!\��2�o7�e�?����a3=�-q�$W�=��)�o+(�T�_n���htgV�I��4�p/�N��hdb���#��P�N�x�1�=������������Fs��bXz�����P_�n�K�_Sg�ꤵ��F�L�Y��t8�{�C�%��F���[��m���8uT'�̧D+=Z��'<ު*�Q�h����:�:x��f�oE�_7�3�F���m�����/��� �T��ܲ����Oc���<��%=0qU�64i�*�.��U��Z���OkRp��ı�c�֟ f��Oq���>L��J|ti��Hi%r@�BM%���q��#�S�e�\���(u�^ �n��>�{G�aVHd�ѻ��ب���Y���������4�=���Я-;������ʯ�M�A+Q��K���n�C���@��բ������J�Qf���I�9K���Ҳ�!.ݬ��ii���� ��.&̀��i�Q���2�%U\��_$m3�%.ޤ�H&��"(CnT�Y|"�}|�+��ÍGP'��S:���|l@�9��}��Oc�9�ٱH�:�g9U7�4�1\0j�.�����1��~����HL:]`��-��r�����h�C� dF��YK�n� �^#&�S~2#�H�@��S
"K�D�x7�FP���9o���혪�7�6?����nqP����@�z�|j��u��Ά$�$ ��˖� 2)#,��ihi�߃=������D�C#t�v�-m���;}UV������d�	*7}�V���@Gu���L�Ф�-Q`�3�PC�.¾�Z_����kU�7P���v�/�?����dYA�:	8����qF���	��`��*l{w+����Ä�ˍX$/�{�3��4Z�K�H���d�>̲%��_y2�TFJ����ͻ�nD�L\�y�%���ѭ�8����0����A�_� I�b�y���Q�Y�-Mu(��U�K�.���@�p�����L���SH���y�s�zg��?v�P!��1���+�PbCJ���B���1ɧ�s4�0�a�)w�w����Aփ�f�g��R������0�ˍ4D6_�+�l��x0�`��cNM���j�Yخ�a9;]���ϩ8j
̈�ݒ�uvD�>���[ίY\K�B�V�Ae-�g�8�A~R�H#���wV	H#��ns*�`�����/P��z25��vU%hUth�ߢ��5��K���@��h�����L�dl���~�F�>n|=�lA���n�""���~� ��٤�?�m�)b��~�r-�krI'��-F��r�z�E2��%[������cfv�֖A�~�kc7v+��-E�[���ܩW�ڶʉH//�-�O]�S��t���3�K"副^�ʣ	8�'�ћ����Y�Gp|�$��-ktڏ1�"���'�8@��aP~�*��p.���
� j�g"߁R%yjŬ�e�D�Q|�j�� AH��~��pA���Ud�2�y�ƕ䢲S�ܠ�W�q��U��}7�v�}�(�R-
/��uu�֠�ӏ�T.��&���uR񮸧5jLG/��<gY[�N��l�[�����p����B�ߍ'����t�t����nF���G��J"*�7�ɲw
�,����s�������ҵ.���2S���p�8�aL=X��^ʚ�*T��v3�u�nrlZz�����}��֊�E �4�3��&�7�6�a�'��hD���� %F��݂WWM+�L��:8	b��a��1�p��t��jL�u�8@����<��D�-����,��\!nCU\g�ˊ���n�����6?;z)G~k3�|R2N�����n�e�lnn��.	 �	����������bIx�zN�J)�l����	�y^�l�Ey]C��(<�׷8��"S|(R��T�c&�{?�eS[n���ԕ_,�E���A�Pޑ����.����(���:4bQܫ&�іp��ƪ�M���St,��e$�3�=��N2�J��[��&� x28K���y+h�roZJeg�{�� ?��+�t�}'�|�]��$���?��8�1���'8�ÿ�S�ڲ�������{����M)��e�m����T�	��i�W�"`���5/�ˎ�rzMGbvD���&��M1�B`�^
P�$̊� {��]�jr�������s魤�qs��Y�j$#Jp�{��~�.F��5�Ȇ�g�q}}/u��Y�3\ՇT��1{e;W�.�<8
)����w�V�P�:�n������G{b@/�1�� K�\.���7�Z�n����ś��8y:���IC^H���b���l��	�A��q���Go��d���=����W%���̬��ɑ���:"*�KY��/���I��.��A�����e��
-�(X&~4A��x�/ ��������I��E�5�IA=ݬu�c糼f�9�F�: �һl�Xv&�3���:�#���>�Jٳ����0���3b,��jg��N���̮e}g�HN:>p��C��Ⴣ]�?��Su�@�f8������̂�' |�^.ڂ~�ci%�����E��/��4��T��ڹ_}�͆���E��"�3J�\�
��&�����~�ř�X'���ZI�	��n���+~Bu����e�VdN���*'�+2.�9��(��󛻭�3��>ތgǦ���Xw�g ����k�F��8�ʤ��S'G�?��7����^���~klؖv�nǢo�I��La���ay�����8,��Rp�þtv�'<כ�B��7H�����D��A��Y{t���KX�2�t�a@���좠�3��� ��ۄ���~���� 3�K22t�䩿�֑������P�5�+��WR��N�*�(Q�O]{'��r�9&턵��i�I  a�J̨���/�O���ͷ)�5=��y:	���GV���G�`����é�WÇ�B6����P�V��4Aۚ^�V���:t�
�f!NO��y9ā��\�>8�̈�Χ
Ħ��DnE�׵1hm��T_򗗯;/�T�`Ķͭ24D>�Q�����S��%�k��
!J���.� ��&W�?�a�{��Sǎ꽠m�5|,��)/�} ����!!\_�i�����&�k�LE�C��Q4S���p(�������u=cg�*���5�@�j�u2��%8_&	'��E���U���������+x�H_�奢\��6f���=����Ow��R�[�`��L�L���������ja����X�0�Gٛ��t�}�����D@�_��~1c����4��w�p��R1�H6�P|9��ŷ9�:����
���2�1�)�vī�ߪ����^'����ö,�������ٻ�r���[sL��o��	��p�\���u��m�iz�<�KՇt`Y^�am�́�NhR$5����R����c�O���T��9Z���5Ȯ^�CqhI�Uh��ǌ&h)s��u|�ڠW���!%�U?'?b�a T��S59?�]�Z"*W�d�'�Z��JG��t����� ]� �t��ny"	��!h��`m�츇��x��N��境4k�,Y�EٺI��ub,;���?	�_�z�Bv��[:^��2K#�}!��X=lބ�����DKP���ڛd/�u����N��1MX�W".D�;A�|��z�z�>OM4��<�Is���,:S�m��e���M��^��Z�������p�4��?��o�2:g�@��QV���!�A���a*�H�EwYLJ*%J�%؅<2�ux�=�0�V����B�k�v-?x�L[��GW��uc8�V��IK?q�U�������>B`��r�o.�����7ސ�tI�[_҄Ž_�,���L%ORi�ut?b!�%xt�� �6��٭P����b喕�X[4:E����k$Mde�F���H�r�-���1M�da7�>#���vL �ی��z�gt����u�f��yc+���!��\[��"�
	�>iQ����H�Zx��LAZR+i� �1�o��S�Z����Az7��h�L�y*�D�}��R2X�$��j�߱�Dx�CN�5���障:��L(H�=���;:�`<3�QOc�,��ju��~d#g=b��E��(1���=���n_ �2�����=&ъ/{��
�v��%�ؓh�r�;���%�7˵��N4Z�H"��o����NB
m�M��` �]GЕ���wV�*�.uwll^5�yih�.���0X��\��9�l�~R�S�^��Kx;�!~$�ˠ⪇~%��9���d\	zT6���s;w,��
��E���#Q�|�f�T%$��v�Ukg�!�7�l����n��cs���g��9K+$�����Z���@F�����}c�����\_P5&o�g׃�מ.�O0�B%��l=�Y��Y�}��/Hݤ���6W������5��� ��5�}��wv"u����$1���J�Y��x��嬽,,�'�®~8��3E��j���{6�����xݻOH0�U����h�m�hjv���Jt��J��J����ĢB?-��q��A@��:i���3ke�ͽ��%���2Bq�pj�*2O9�QJ��@��!����f;@�֞��̮$���d7�Ӵ�\UZq��$����.�PP��_+,h0�SH��8Mq[TG"��l� ���}�nvW�5�������=�8���($���[�3��\4#�}e���Vf�f\�MR�{qx@�Hb6M��
kK��E���Bbg������h0�MŬ'W�N�'f l�C����y7�(�ÇW�)�5&��X��(�Y[�l� ��f��脲�L����Z~~\�}����m#���73ܼ�� �z6����.`����zC��;�4"��"�@�S�U�h����T���2�aJ3�hX�D|����bWh�I�;�V��-�J
���p�Y8K�ŏ��[��>h	"�{&(�͆JD I�6�[|��]��C6]I�h�[�y�"�J��������]b���o,=��d�ֻ�Nm1�u�n�9���mv��W�T��Ϸ��~�5_�7)���X��!ښ	@��a����J�N������u7L�v�s!Cy<E���QƮ!��֪�|�׬�/6�2Z�J�<�E�i��	�)��d ��i��^��LIj�>��AD7:�ۣ�o��M�p+G.��>����P	ShrЛ�J0�[j���ʢ]~���ZMa��A
�=���A3�E��F�S��yS3��*z5�K��������^�e��7:��N���:�J?L���f$m��a!�.z1����G��{�X��r�=�N�t���	~�ޓ9d��;:E�;������WJ�h������:0�����Z�]�`���Q��^�m��yr�1��&L9���.K�Бu73A`c��'�
�\�d��AE�>M@���2i^5tʜS���+t���w�R?2�&��2h�����N"na�xEd7�����bH"�'s��.2K*�2'��������[~+��׋ًk�#�\I=�����wj}b���azv���A)�Z���ď��}������Ȥ���U������Lkٳ�L���.}L���%�E�c{��}qI?�?>2���"�TG��Ql4/�0���ԅcz'hesMrQ�j�9G ~��-Ҷ��<ψ�xc"�7���-���LK+|����~У��Tg�� ��_�ȕ��ֶoR�n�OдŚhy)�h���i�%xd�L<cs����G7NsTf�r��	�r�H�7��(��h�unbHly3:��&��^g����F]R;eP�1�Ƅ�ݞ�@<�s�p�o�ȫ��*a�~/�������r����2U2�I � U�C=�*�X%�����p{,\�4
6淍w����k��a�6D���pU�( �������h��Jn�1u��}�"Q�����YAd��P �������{/�/�0���no���ޘ���6�2��9���ɧFV�����=]����~��cS��&EP�z�"a$@�{�E1(/%�N��6)�<8�e�k��=���Bï�}A��8��}0����ڪ��E����]��԰v�����9�PbE�ڵ����}�.jL:�ςu���Å_�=�q�@m�^���g�m`�-�qS�k��:�D v����`�T?G:;����sDn�(3�� 2(2i4{n���,�nL���^�^&%����O�a�1plE�֤�wޗ��	�g&-��t!U������_���"Qn4���O�U�!�,�-��T���s�ug&�en�vCR���I�0(�}A;��"/�#���{��%n�������!�Ud0������t�B@��f�����<�F��Y��%Gn����?ŀ�$畣aӄ�W���ȇ���������K3����}�ĸ���M����̍��\oB�cn�겾P�e���|���<͂8�	 ����UON��\h���$���(Y;������Ʀ^+ҫ�J������<�Q��Z��,5"�]�萼X"-�ދ|컼��f@Y|��H�i���<�x�wy�끑@�&t��q�-ټ�~6�[�O3���<V��	 �K۪�W�/��_�'�O�K��A�|�ė���qe�A����Q��"��"���=\v�q�a�FI�t��S��g�!(H�|C������+��d]����4-�9m5������Vq�s�Ʌ�1�l�?�{G��Bj0M(�hh{[���� �5W3Pӓ�Y~��"1��j\%��.=��1%��.� �ղN�5���2NK>BdxS�=&��A�(L�z,u��gb�n)!Y"4��S��<������
 ��IoZ�Ҍ;�Σ݆��r�m�ΔP����T��m'�����D|���lDj��R3���k�j2��$����ro�ĎS��pO�i������2?���\������L���Q8��vt��i-��i��e92j�;�0h{�攍����1
��L��O�p�pA�����J�}�^������ŉ��.��4\��y"j��Htw]����fr�_����Ї�N$M��ܦh�T��\�ۣ��nպ�q�'F�����d#9w��t^:�䇖�$y�mq�8S���z��eq�ɟ����@�م��+��dM�"��Չ$P���{Zh�#V����p����K�7 ;��FKq�u-����d@;&�Z��;W�$@]v�!\g�����Ҭ���E��l�vazMJ0ix�vl�U2����3�H�گGL������r��.u�z��֙d���,�` θxg��e׿����	|�ϧz�pĝ�-�GU�a� ���
萡3 3;�1�i.Rt�Vt��-���HM�'�*aT�!�^B�u��G#���?��ꮛn��j�'f�G?_����m$���$�k���6��"R��xzRg�*�L�s*�߫�Y:�O:�����:�:����`���N�	��~m����/�=�U"��J�"a9���\{�����\كA���
.{��s<�����/r�W���	�g�:�8X�Ӵn����N����Q'L���}*I���)��Դ�'6b���Lvxy��-B	Ǭ��16a6f��G��>,ɎL��BG��u�q�<J�s�A�R߁$��W�����s���Ҏ7�VH��`��D���,��+�^��M��p$vFTuo{�� ��h[��E�]�k�g�W��(�h�z,�V��~�>��p�K�z/0��*XV����1b��xR�[/�,�x��4��%��b��px�JL���Aڑ9HJ�k5�Rq���偓=�п?��%~Fڰk!֮�N� i�2o&��pm��v#L���Ո^�,t��\��R�#�_h�_��d�{�I�{�1���i� �r�qp��UU�q7�Hޫ�����T�_�NYH�Պ�9Ln�`�0�Z)�uz� �UTS��(�^�4§&���v@S�uI����[+ �����M���ݘ#�u���M� ��:��Qx3��st�7cy4�um�4
�-�$M�\�`m���Xl�vi�mnG��/ �Q$P����{�|$W�&����ߥ��8���Y�>���G�
�K�n h�
o�g�f�Q�Lw$�6m�=��ҏ�(?�m�]��q��g��~D��5��)���UN�������c�YX��|��*�w���CAXF��<s0eLڦ8���_�K���2c'ROF�<�� ��j��Ρ��`��)���ty,�ؙ�:�N����)���H��{� ��O`����FVr����\,���s��!a�|
���5�@'��T�{"�I���
�P��H���?���(�����c�Cɦ�Ȏ�Kd�ܖꢠ�-�A�F�<���Gpd{U�
i�?�H���9�&߳Ⱥ�PJb3,HB������v��d�V��}eiW(��!�)���6;�	Mo���$Ĕ E�=篆Y��[3:sg?�a�¯�̱�D��sJ܎��헋d�f��F���A�)�2ё&vg�|o��Sԩ�M$Z�Ў�N�X���I��X��.��3�)WO��b�^�"�4�U�� ��Z�t3�$w��@��&�,r)�l��{��b����A�{��n�A!`QQm${0�ݘ7�O���%��Â��*�5�C&�'/xP�z���-!�مI�G�����$yUpA.��4I_�Y�p��2��v��i�T��USZ���ad�P0���/�(R��_Z��Rm��d�5Q�I��o�љ��t��80�.]�w�� �d��1Dd��3�\s�IT!� �y�zBMG� ��/?L%��`7���hʧ�0u��GjS�����12Y6�äO�*���SW-&�w�&j;�����f�JB
ψ'Z_�a�~��y��κJ��VA� >�ON��_�^��:��� �1���k��1E.a6I7�}���d�M�]��k�J����Y��"��R@=$�9��l�^-���l�Õ�����dJ�a�(k�\����}m���:�$b�W��@itaG�S�(��&��r����CX�����qy����>'Sb�JGf1��|z��w7���%�G�^��	�s�p*q�A5h�=�H@np~ �i�l�x1��H���T�Y~��nPT�?�s�gb��'�`�������T�kU|h����@�R	2m c��r��4oJ6�D!�We]�W/]7��#�8���8ғ��_z-}�AY�mm����W@��^�k��Ouw�\������)�sq�����| xI�̿-�Ț!҆y�݀��.a�k�[tK=�����2���|2eE���jak_�*�ՎM�����~+nz���!R	����X���x�I*37wTUZm	���:F1���q�_���e���Ԥ^��|	"�un�a6	��ǀK�Q�K�M<��ї ��v�����e�{��G䮀S�d�������Wv��p�U�l��KMl5�v�赬Id�(z_��A'�� 
K߉������tKx�(\��	��.�(���P�yf%mᘯ���=�eP��&�v�h�ƠO�#oimOfu�j(W�k�_\8��醖 2+��Y�^�6���ď���OI<s�L���PɘYF�{_���o=%���E gG;u����8}�B��$8���H9��TL��?���w"Ի�N��s�B�Q��l&�qn�~�FL����&}�~�z��`w���p�U�R����5a*K�	��QL=���X�Y2
J�:f�����?�i!�k�a��.�O* �މ;��l�K%��+?� ߳�*��EE���
�M���"Jd��eZA���a�=��'�8W"��C̠�S�>;��tF�_�`��Dn�M�(Q�U���Iz`�u����`=�W4f�5��3����t4圖5@w��U�oq���i�D{@7{T�����ŮF9	z���Tʋ-P�&�f�@�p���>(�8i�^��O<� �	ϩ���4Pz5R�;�������iyz/r�4�x�n�Xd�Cq�T�V���1*��ƍ��6�1#������ts���`�(��qs<U�F�_�L�I
�����=/mz���~`�.7@�O$�M��0Z�h\��/$F�W?$�Dd�&w�uɟ%��f�qix�*��s�D�R��h���W߼�h�����K�
Zp�WGo����m��_,��k4�̘�0�f5���?��ʹҵ�rj�%�-��g��ۋ��'�N
�No�0S
�[�"��(5".� �h�|{<	z�wqs��^�	=tgmm�yiS+p\,���A`Ӵ���fg)���AV���Yd�Edc���,��O��ّ��=<�0��1:�T~��3�����(ĳ�3�0�'��������X��g�V�s)�gU��6��0�'�}Qd��e�}�x�Kv�;���G�jĻÓ�6��a���v��?�'E������$��`�uB#;�VFM�e��E��g\��,Q��$m��t}
�n%,5�a_��p���1K�
���Eo@�q�WA�1����B�tP'�x����`�Z)�gɝ��l�h���1'��V@p<uz�cT�]�|�������&�n���[�%�ֿ�RմPL��N� �'^�i�lf�����Np�ƎZ2�L���z�=VMŀ�9��4͂;S~����Y���!�͎�䃫�	yt1�"�B�T\�kW����q��+�|n�r��^��\��#�I|�l\�:.E?7X�*�F���Ƥd'е�[�ƽS��7��M}�y��H��S���<F�{]A�5ȑ'\�v�˩���a�*f=�j�N.� ��i���P��4��: �vU�%HfPl�R�5U�b���P�4oc��[ �g��a/����!���H�a+!�q	��O`8E�@��*�[���x��ਓ)X�4����+� j���N*s��b0������KN}�
��	(!V�;T0U���{�;���T�&����v��0���yW�[�ؕ��J��@$�d+�;��Ml�2��H ����]�qzl�ڍ����v�-O�QѨ���O7,sf�����;F�,�
~=mbi������Ș�fv�W!G�ߏE��뉓�uh|w�p�8��8��]�2��i�S!u������!Uә�g�
��#���PmH|�q xv"_L�Ɛ �i��]n�ٳ �H!�- �ȍ{M;po�ć�m��H%H�>��k�aw���t��0��?�ô��w,��z��Hg���&w&�w�쪠�X�"�!'%�:媨��gK��e%�8jV �#�,dy�@��%��m�{A�2��%��}�ڴ|@O�a�t���b~[��kzlUKa��M3{�Ew\�X�H��滛XG�O`B���F�p=��=h�J�y�<@|g�S��� ���d۹�b{\`]1�(�E��E]
7Vz�˱�`"��p�R�Xӛx���*�։G���7��j{��Ͻ��݊&��M�p�P���K!s)D�2�~)n*���B�(�tЕ$�☎1���}��{mq?߿�����Y{�z?���<{���J�q��
$��1��{�ا3��c���p٭0�-"��Ŝ<nd�*�
���n&��â���һ�q�J'I�D��[��r�+���<+�2���y�q�,��IK9�}v0;H�j�x/���ke���a<�@T�ǀ4t����H���Dl�ytA�F����i��K�_���n���
��v��<��<w�f�	�K-��c^�:3s�e>O�-J��@}���#僀�"Yݫ�W��i}#�,]�w#y���CO cU��l)�=/"����Z#�KRh��=nS#�Kg���Hg�n�����.JA�|ow`F��)��X�$a�%������Y��Lqe������a�T;�7���+����s��}�� LC���x��Tpj���)ɸ.L �Dc篽��b(�9JѶ�l�,J@�`���d�3vx��XW�0�����6�)��?�ꝱ�d�e�D�in�X^W�e��.p�z��Y>nzs ZM6�3��(8-Hϭ���-�˗�^��ܞ��$���Ci�zLa���Gk�����6ؔ�p��:m9*R_�ÿ]4G���$��mH͌۞����E�����Od�:�݄BI��*~r��[�B��Uc��?��!���ͷ�㸻^{"-�{��y��=7]��vM�l�������H�5��B�&�i�{��+}���'͆ߖ���X�Q^u���wv�䀯>Gm�l�.�������	�b��
�D'����:�3�[��`!����6�BU�n��b��B2 �!&I�I�T5�����М�?;~F�.}�ߥ�]��ťKr���-Ǜm����O�Q��t��7�����|�.Aݟ�X�<M:6�����j�3����F��+�+a&���5�d^=��~����~����~����~����_��px���2q�}z붡*�v��Nyz`�q/�R��'�TBJcz��nX.љ���e�BP���Mѧޭ����;]P_��Ks�nr5�r�T��!T�#��6U(\߾�\�;�r�o��S_Lԩ��_D�NX�>�~�#�F��1�+���W�e�.^��{}��tW��$�����i���E��7�s7R��M6���tä�Ͳ[��6{��:��ft�w��:)��me��O�ʋ3�Z�b٤�I�2���s	���!��]�	��L~�tdge�r4���}���|��ir��c���ϥi�!\�#������R�!{X�+KZ�-"��"|�O!Uo�NWN���+�5$�Vۧ��)�X������zݙP4�Ċ�՟���&z���I�����o�L
�N��6��1���뢻NyV��|�݌��\D�#i�����Â
�4��������7j�|#�`�(U�����TS�8��,+�	p����^��j��Mf:K�s�"*O��{�\�����,�lN.ڻ2�����17����U	3-��t�ͰuD��W!~q{T�b]�8}��t��8�Sy��y[p��;H��7�?ZڛHL}�{e�j:f:�a����c6`p!/ $�꤆lBf�\�b&՛�#I�.�N�h�+;얞a+$�۱�t7�������6�;�kxW��y*��
m��Vb�:_N�KԌ%���Va� ;�輀�y$YՖv��5���~9��q������&�g�>K�DJ����\y��F�<ƃ�w �|�r�����y��b)3<?G�� �H��K���y�Պ��Z��'@_�]����KcKB_a���-��Ѷ6»�]��0e���I_��d�l��q�lr>q��Y0��4�b@�f�m�Y������w0�.���f�,(��A5�z��jK�Js�؇2M|�m��H��Y�p�N&Q�������Dn�����[��z<��h���URr��J#�ave��6��u���S��V"�s9WR�隆�,���w)�J��nA�_�N�����͎��/���L��_1`�P�o�z�$x�JZ���#;_*����)�M^[��ۄQ��=��ApO���쭔�K9Cv�~#����=�1�BhJ�w��P��>�F�cv��)�Q�fD,�[�ˣw2賾=��8!�G�5q)k�J�d���:
���K3uw���gjD&�Y*��}��G����U.����ml�0nM���\$��_~Mz�M�o�z_�w-Z��Z�Wp�y��>�9����vY]�����W��sS�N�o2_P
�_*�]g� d��s��(���&,�qn~��a/��kZ'�J�{�N43	����l��n�o���'���φ�f!̓�m 7�X�±��ey���p8���Q��?��<({&T$���� �h�ؔx��b�d6F+�f����v��S�[r-��wa [�Of9�����wN5���vg��C�}h��i�����
?��;�I�6��S\y��
fǿ��$��٬\'[�,>e?@��ƣ?v������	i-����6�Prכ`����f�ݜ2'։���l�!�*
/d��'���ü�*����o4)�vQy�+C��)ߡ��TV!�yҊ#񊆖2��g=��̚��٥�	��N�mj�}S�� |�F� �G��n�_��0h6v7n� ��=4-?�\���������!�]K��Y|�hK��ڱXo��}oBr)5���ƪt�y6�&��et��!X�Bb�aB�?}�����~Ո����k�7^��t��ƲF��K�7Ȁ����fEF��ü0-�!��f�8.���GT��y�$U��Z�3����	�?'��4��q�P�2��̬�jtG�Q�f+c�gt8b���*H-�t���:�7���� נ!t���04��iĵL�b�s=!�@i���ŗ������>�/񆀝?,:p�l��49����Q�Ox`���;��MzR��HP�q~�����ּ��>n
d����š�N�1�v���V�2�ޱ1�`�(>[��Є��Npth��̈́X��8zTC���H���:��A�U��p����UR{�K֘�J���o���s���}��c�p���6r��b��3:�κ"cYO�W<�(�L��;��l���p��o����l�$��	W�\��l|�!ܩd?�pK����
�&=��P�-�� �>�+��Y����� hS�쀩�_�:�_�CrH�n����=��T_����Y�/ޛd��U�O�X9%�o�]f��j�*�ņBv�F�0�ԧ��R`�q�ޖ��`߲	�J(#
[�%�_�<����I�Y��g9�-�ߌ2Z�
BU1��hX��D��3�@δ�r�-�UK��ENX��0�Id���H=��4R�Md���k�z�>������->%��OX	7Z��˘
��jCH�խ��OG����d.bO�,⣢A+�v�9��������~���C%�����~-��D�T*�+��߸3f��K!�s�p��3�a8�d���mg�<�~H���Jan�R���B����f7�eL}8��k��8O $P�>Ռ�A��#sH���1N��'vK��ӣl��g(�Ω�Q�:�z�g�%6�@��'�^�_���Ϭڈ�M��~�
��߲��!��A�F������q��r�盆F�;�������(��ƒ���28��
~t�rĞ�Me�qE ��U�p�s��a)��jԓզe5¾ g�!�N�������_ٲ�݉:X3�?�a��V����5���l��.��.���c��7����a��������c�������-��; IFL�`L�Ӆ �[�]��jG��AL��C�������A��Sn�k�j��~ϐ��Hl'�����ֿ�{
�:�[j\g�fHDcfn�_�ڴr��|��yOihً���f^��&q��\B�J�~f������s�KV�e���:�>�$��i�_��j=Wr����s��Zr�g�U}�y��0�Ya$v��nw��F����Y2�Z$=!dyJ0��=Pk��p�d	����{|Ӛ�z��@A���~#,���EP���rR�=��N�E{�N��jH�N�;�LC��{b��^ӣ���~g� �)#���A����䐱C�G�EnN�?�n�q�2ع e E���*}�!�a`�;eņ4�	�Lj�2�_9rǸ>�y�XX���I�:�` P�[���grea
����!����s
�W	��Ѹke*�Ϭs�u_�7Q��������64#��Uշ�Dt-�p��M�ټ�@��\k��50j��
��l��1��c�ֹ]&�ES��x�.#w�
W<YQ{$�����Ƥg>�`��������ެ
O"2��|�%�fb��q�� �U�{���z�%t�j틬�0q����1s���9�aZ����ELT��A��:/�B�����A�k�b+���0���'(�)�
��B�-�ʡ�#�^/�'�c;ˬ�Z@����qc����?	Sߎ�f�# �b�0鏅��Ÿ�kZ��G�P��3���˙@f4���@�09�� <&�m��S�N4ƃ�+���}�V��Cd0Ea�$wVq%d���tD�ѳBH����)*�H��e_z�-s�`	F�=�9	��7[*)wx_�=:��������P5L��Ty\_�C`Y��dIQ�emn����Ä��0�/�/�
Ku�D��=�����1z{.
�Kt׃�㮳�vN[!,G�yˆ�*���oS|�j�\@�1�wY� M�g���qyM�7��j���K�\r�́�n'VY�1�@����������*n��Y�f�x���P~�%�$ż���DJ�/O�1�^�I�ǜk/{��-�ÜE��Gf:\�i��M�������؇��$���?�|�w*�Q9���v1\���S2�6�G@za�
h5~6����d+�K,�·��m�ue��Tr���>���c@^	�j���
H���^+N_�E���B["3�-�.t͜��s�-���̧������~�e�'�_�=��{�U��g��s��Ѷ�������Rm���^V5X��MwI~,���B"_�
���<�O���d��T��S5os��9�͹�|�ٌ!��	nS��Z�g͡r���L��s���>��1�? t�����JP��Yx�I�ؐ.�$�i�1|[�~N:�|R�̰�C�o𮼃��r����U�]����SԹaӲiI��0(Y�I���I�xM��k��AX��B�8w�:�P�!���m���&1�g�2������&��'���$N�q��4_�4��mH��b[k}���`�a ~vW��ML�ďmX��O>&�.M�rV���"?8-55��9�����Dg�o^XY��wL���j#�m�I��r��ei��e��$��P��%�i������t`�]9�!��>N1�����;�	@_#��Z�S��3����/%g�]�76~�mH֯J�ͨn�
�A)J�?���K;�.�/�+P�YseА}f�7~Iu�FF���sM���6��6���/��s_J%��*���JͰ(~7�����ݦ�KYA�ν���jfg�m�&�׿1��g��$���1������v���0vD�$9"��xPtp�T�Ю���R�(d e1�{ZE����&/@P�Шs�
g���5�G��3��j��VA��"Ĕ��7�����
��h��m]r��
���8{+}��Kǥq|�P>�5Q�j\�oxg���~)����H��$�*����L�?��<踫��2<.�2�HZ��Eȧ� c��oKOQ�����6���,snq��i��,6��LB@��5Z�`dh���oC�`B�����p�ar�6E�ۋW$���a�^��3s���ҜS�5��{d�CǾ�v�bq�f���e5�����b� �VW��\��3�������]�'���m����Dq�1�~X�3���� �Q�����%5u,��'��p�B'�\��ҥU1w)L��B+�2rL��'��z񷁻8Ƽ�S���4���tpaUe3 �|��~c�0!�����Xna���N�^d7�)��YߘɅ!��S��`��ШԿ�E>$�n�O���mGmM�4w���N2;�X����W+{64�8���䦲��-�r��� $���x�4�laH�FW�7b��'D���s�0��g����s��=��� н�6L��
��	 �:��r�%	�2��رA� �Y�:�Gg��x&�Q�<Q��vxX�ȿm|������H�FKZ�1S���N:A�8�H^�-G'�kDHaxivq�Bm��[)>��Z �2��t��G�nK��J-L�.�z�/�7g��s��B�S��,�W]�[^��.
-�t�ӵ��>ʨ��!)1%�;�o���!F��[wu�<�B�y��^K�X���J����P^#6��7H߃{���?�+���E�垫�]�,Ow��\���n��(�,�\P��n���}���s�sВ��/�ث�/䠙�G��+�"��$����oח���$�s��V�v:�$��x3|�v�3"��v��@GLj����:0p����S�w�lA��@i�y6q�1M.�$�|�a����x($�k[z�&d[ۃ9q��.�V��xw��v��E$��/NT[��V̀+ȝ͙�L,��ݦ�wbXS�'gf��rE�Ca�>��vbr��>��b�k�RV#��Dئ�Ѝ�ݪL���(X����6��Iջa���u�x�S���k�'�*C��3�3�T%��U�����'V������(��0�]��f����΀U��#`9<#zS;?W^�yP�QF���<kMG>�zV�]��nw��_.��z�����Q8�����X���}{�H� �1%�[{�p+��0�_NrSq���U8�.E�*L��]+�qJ�Ң-��#��;�JV��@S�%O�ʻm��k�)�$����"Ķ��$[U*Qm��U�Z��"tJB�H���c��Z�=���Hà�8���<�u#��~���~(�|�����),r�:�=%4�5�F~���"�Ũ���P�r�iq�[��`@Qőr�o��J� o����Ҥ���_�Wf$���*8�[Ė%MMК����m��?������9�M��'h��#���pfZ��%k�Vn�a�G}ʲ�3��"���z3�~~H6:Pv�Z0�3����H,�д�|�&�=}}T����!�A��kб´�%g���Uom�Z��W=Y�a��c[�xTR���V��w�~���fm�&�p�����n"�������@��2-�F���_O!���J�[��`�Mj/ �^�W�������=�	����v�oq!-G�ݗV7�9�h9T��y�9Uٵy�!L��L����#QV�,ceS�V�}�~$���]�z&
��R"V��gb���l~�3�hv;�z��5w�o�e�ҿ��1-�<'�?����t�ݪ,��*x���Q�Z���1�Kpjÿ`H漂�+eeW�#�rC��+�ĤYi� ���S$�=��W���;���
i�ϑH}6�E��>h$b�w^ۈ�gg<�PR�m)BKo��?9���1�-�9.��A���MQm��M��x:;��ib���ͳ$�R�	�X}��Ԕw�M���*�;�=�;��� �Њ�ڊ	[y{h �*w���i\	�(U�hX�&s��b�Yn��$�0�'U�,j�뿈��`�,2Im)��ƈ����&є{���%��5Y)����E� ц��Lɵ�!2$3����M�W�A�;�x�fG��#��8��^�e�/�~��~��&���r�1��+���T�ѭ#��mm�q�Fb-A�MDҢ��������9�ߙm4���"Ϻ��# ��Ru�E�0����O!�%5ǵ5���ZiV�*ň���Ji�/����Gz� �Q:��۷W�̈66'�������hZN�l8b�m#(�f���O� ��\0�����w���4qVۈZ�&�/Pl�6h�F�|��U`�'�&��h��Vs�U�������H�_�66����1&���D7�ma��8(��'Am����`�|��L`����ᜪZ�؈�m��֖I�d�r���!��`���u��WҐ����x�E��$R���p�4�$��dKl���m�\]jO�5��^Y�$%�!�?���3[�B�v�r�֪0ls�N˥r����Dp<����Fù`큒�F���+��8R�S�0W*,ah����-bN?�龥M��h욢��7j}�(���wv5�^1��$ x�PK�y�E����vX3�l������,�%� DY�;ąj��Gߢi��X�O�[Ғ�[�U��T�KX���5�x��s���wf&کh���-�^[�EY�ϟ���w��H��ȓe���=�|��
c8	��^[n���,�#�e�"�s�-1,L��;I�M��ͭ$���b"ZAQ�"ʤY���U�N�G����-h��3�F|�J�l�*��Iq�$!��4B�Z~�Vp���nƴ��
�z�N��UԨ�3��T�LHq��ʈjW i�GX�����$?�'�V���{�S r�C-;[���+3J-G���7����#�.F3\��c�6]��ӥU�"��C{�G�U�����ch損�׊��3������-[���0z�a<�=�x9C����"|�ȼ���]�n����)²d���$I�HbT՟\�칔Uo	A��̳<��0Aq"��D�o��~�5� \�Ÿ��Z��6T�����羆jp�旅��Iڴc܆���Ί�+�lfب�Mjm��DOz�n�6[���hmdI���=�֤�䌻+�3k�?��v��pr�����+=��k�،!ѓ�|��B�-� l�F���[���(\a5��n��^;�I�*1�,5�ܱ�/���2Ȇ(6�W��j�ˎ/���ҵ��:1�Ck������l�w6�s�g=Uϸ⡇gL��&&�f힮$��~�>����@9��J�D�H��������`M��*�+u�'߬�WX �%�3)=o�*"���'0�$�q̿��$���u����'}�!�����&��z���C���/��
�O?��?^�p��ɕ9r��S�8(*H�� ���|2Կ�}^���	�(Q�H;�R�BGZ�ù���hD,q��T1�S{�{�-h�=2�"j���F�J�t�ƿ�����Tv^���m�Quf1j�/>����YGN�}��zw�|�m_w�����@���q��I�qF ��'z���HǴp�"��H��O��B�1{�!�oX��`��k�C��v�8^Jpa��vs;�q�!󖄡�#����S�� �����!�, v�.�'�R�}Md���Lm$�F!'�Q ����j���
�z��2D�ȏ�n��Ӣ�m����ȩ�Jr��;;8��Mh�n@�%v����N�]��' ��9C���mb�q��o�t�h3v�=�.7K�?��5�U٬+G�O!y���P����2���V�!
��?�)fVQ�pÚL'
��}�x�6"��\�,��+!��9�+�|���Qe���X?m����Ϛ0�T�"��JGd��5�k���k�gD8�����{�$�3t4K�	����ؠ_��F��y '������_����3i�x����Rg$����{��oo��ˁ�˒��.�@����X���K��^��\�]V�=��ȫG��\Wj��_�k���RS#������H{�/X�"�i���a\��.$��|��0Kj �L���~�-�ЇLRY?=�X�}p�,� ���Gxwd��|a�$g��I���J٬��@�Gʦ���ė���Fi�5ZA�J��@��ܞ�Vȴ��VFL��Zy�6 9���}u�-���5߁����P5��T_%�;=���,y�?8R�Dc!w��1���~L�H�d\	�D6&-�K��zj����_ �,&�X{.��,�Ď@vZU�;�.�j��t��~��dᦁq"�m��_1u�4���Y�����/���n��h�ߓp�(~���w��v��rg�,��F�K4��#`����=4o'
��X^��c�eh��L�E��q(����UT��PVx��˶!�MsZ0�Z��n-� ���|��[�-i�B�2�3�����J���ڂQ���������l���2�~�$M`R�b�A�}z%%6�uv�����џ@�=8�1
Z-n-�Jm���m�+��NF_DKv��֬@HUk�`6�g�ԟ`���������2�aU�bU��ki�؄�$��3r;�x8!� 1�em��N>!3����0J!%s��uY�2������Y�n7X
�M�tw_�"�y<
���(k߲���+и+L=�3	U�ކ(KZ}U�����V��J�}�d�D\���U��= �>^��Ô�;e��!@:�\ukjm�I���v��d��7�Ģ%g��Pk������7�:͍@��_�p�����v�F����y�;:�^U
Y_�,��~��3b�~�T*��̒bt���U�@Ū@IT6ɜU�|��:)N����[������σ�V���F�:	�&h��V�K��=�2xP�x~h��'��dp��b��G�vr�z#�����SۅA�Bŗadא#����+���{b����rv;���'X�}��o{��E��7�$�"��Ɗ���q�׫��c�+^��|T#����(d��ѓQS,i�8��-��OJ`�����pW��ŮM�#MK��P�VX���s@�B�6䭵 ����_����|���[�$''d�-� G� -.����G� ���� �ʳ$24��_�Q�pX��c5�N��a�c5܈��_(�F�>n9ܤ�c�
����FǏ���Ӽ�^���}�|���y��[/_�29�O��$��o/�����m�Y���C7�$����9R�h��<+�>���~����4z�c�5#�ޑ�m?�Y����z��i6�ߴ$���-���3Xz��r�dd%,Ǉ����'���������vD���.�Z�hWuلg���0��o������Mq�Za]�?�yc9��k�rK��Mm�G���b	��l����\���l��l�U����7�Wr����(�SU�`��<r�y���/K����5�h�.�/ff��bĨڢ7�<���Q�@�6E����f�ȳK�"�0���f?�\���7]4����rX���JC�f��z�a|����9\� -�����R��9ߊ|]�M�l�v�D�C��N=NUB���<�DG�`Ǜ�s��H:z�2By���Q��҃�p~�+9�;3�[��ɢ���]=���I��-�x�8"1����o�ɛ�ؿ�~ɧ��%]�0�����ؚخ�_���%������P���PW���hƪ.iR!C�?mS����U��dئt�%�¦כ�c�	ǲ)��`�)�ft��&��UԤ���[�:&��8��p�	G�RR�NQ���.O� �ňİ	^�)��x�9�տ�7GȲ|=q��Σ{l�?ߋ�P?�~Zy����D�yW>�%S�߈3H0ݦy>�r�,qna���L��o���K���g�$ݘ_o�����Y86s3�W�̀�ǫ+�ON
@�o{��)^�D�/���;Z:~c<�[�\�3m�ݦ�����ً�r���Z�w\آ@��H�G��>́X�_p��a�X��羅󆖌`�l���ֱS_4f�ޮp�������'��j��i�F���y_{����1W��E}�%�r�5N�s������Ʃ��?��x�P?�~���C�t6��+��m궳��5�.�~5�є9SR��.ǌJ<�0��{۾��Ӕ�+�X��.G�>;��V4vT���+@�gL�*ϛ`��������7eC3U��=b����k���~��/	�_;�1,?1�(����6#�.U�v����W-N�X�V��k��xy�?5W��~s�~m�9����Ei��~�D�V�I�?��m��saf���(��#w�B�v�LK��|���8��UTL��k"�iރ��P�w�������T0�	�1��G�JFxb�)����o;�[}rd�ޢ�H��~�)2��/�?��i��Aq��W�١��C�{)c`��������ץ���������!�Y�ȯ�Oh{M�����*��n�8��'���xg�H_I�ȈP~�_[(�׮.G����ZǶs��Dψ.^Tp��S�U}ԭ�-k!\}��J����[ژFy>dn~��/�+�������p!�.��>n���ӓM�����h�O�W+�
z��M�~�em�d���f��ی���d+q�ɧ�[8ˇﻄ6K��P��7�p��i��l����F��6��ԕ���y��Ŏb����?:[~A�V�2#'?��W��k4ص��QZ���]�h�?��
>�ox>��l��-S�G%T}���ٰT��Ѱ��ی�=g����N�y�g��M�َ6�e'���ǰ�G����δz�J�zW��ޭ<����(|�6�-܌`ö�o������]�y��ٮ�@��M��,5͛�L�������/�]�������l��[#dC���O��Wg�P8��~G(�����Pq��[J#�|�c�if�ٲ���y6�U����Y�o���W�6��ƛ^ ��N�Ʊ���O��=˃
[�-�Gz�DU�'o��m�����q�f��횫6��w��!6������L��n[����0�җW�t8��B�?�l�6R>]�ӂk��`TNX���G���Tg[dr��*�?��y��xU���z���5�^�����_�dO������ĕLe��>̊x�yâH��t���=z�)�;��o�T9v����7.�Ai�~�)��\I�~�����|^=�=��l��yMZBG�kr&2��oz��A^�_�^�7r��z���װF�y�0?A�1Yɰ
�1y� �3�bv(8�I��d���\\�ͬe?����TF��a3���.�A��&1�
m�����P�U��/�ӉV�D�O����R�g�Lv��F5���=�i#�Ed��s�Ea \	�����[4��X��G���T��pБ2�)@�|�2��S$��6 ��wI���E�v����I�
!������n�����߃wX�Tt���U�-��]!�(��Ě5%�/�v�J)R�S��gPשQ��FA*|��!��(`9��=�.v�vh�xM�XoVx���34��-h̦����ǎ�	��4�~u춇ƌP�%d��������3{_n��t�M�ă(Y�e���x˗h�j���M`�o�h�ss͹>��PaR�)w������qN����Vg�4�Lt�(���s��=�y�{ �x��,\zlŹ�ٗXo!�T���k��F��jZ���,h�<_Y�Klz���P�|�o��GlU:{��-W���P�I���r;;�M���j/�"2����*eo��٥��(å�c�%;�h�5:�(Y�8�Ő�ښQ3{�~�����5�4	����I���a���Äw0���g�;�&��NƄ��=�z7�n����M�&�հ�>��T�O�-@r>}��{�ы�촡�w�5x�JcU»��ln8Ě_䀭4}���5<����=Ĕoa��w�ң�H����~u 巫�?Dw���P��e�%�����ONyﳕr�Q���YY�96�3��`��%je��OM��^j��<B���D����q��LS��5�5H3�n"�����F�*?�KU��l�P��eM�"y+������G~��</?em2peU?Mf�ZEs�8r<*�u�z����<�� p���h[(���ϟy�%+!�㢇|�����<)=����ss�&@�����E[��`W]�����ro�+��H9������a=U���(l����'.��۸9��e����o>yB0(t��L�����+���U�����*��␍�
/U�1�E{����h��wBygT�MU����@��~���bM:������z������c�a��Ѹ����n�T �\ny��Sh]���'��)z��n�F�s��8���^�eg���v
]1E�yd|n�m<2��T�f��������1HB;ꊐ(��#Ӝ������c�������N�-g��n췼9BN*�#?�7A��������R=hE3�C��:�ˑԊ�&˪@��p��/��0��htyJ�#�˹�v
i#8[�xs`ҍJpO�OD�A�r�aF��S�Q�X��ks����:�`a�Z-��G�;_J�!�|���R�vNi��rӄ�~l��L��4�$�5T	�ԅ�1��%��6pb}UF���Ȭ��������� x9 C����<�a����]�^-ݜjr'�Ǚ�w��9z@�@.>v1�4�,'��K��h�L�i@�\ S5�� ����p�i�6��@�E�]q�Y'���XrO����b�����I����./�8[o4�s���w��<�LG'�Q� �H�<��xPprQ��DJw�	>9��۹R!-;�$ h�l�ǿ�w̢qz�;dYJ�Û�������C}yHdʯ�6�/��/�|�w"�lC��u7M���^�!Q�o+�l���B�e�P?�ʺ"DS��x8)�$��mǳ@Ea ��
d8Ȳ���8e�� g���zrɂF�<U<ւ����D!��w|7��L��x=5D�^��F�m2�@ǂZ�6������}* ѕ�5u��_��}4\�����#Z5���F[��/�ʼ�ܽ`ȍ��FS1gl)ȝ�ʛ[@\e�[V�(ڠ��hZ�@�t��i��@&ai;yS�dd�� ��NY�(��к[�xW��c�s��3:��H���]���_{kV֌��"�~vf�%��Ȁ��ۻ���\�_�p�w��5;�t��^�����G�}�� u'�z
s3�h�?,M���)-�T��Yg�P���֝�E�`C�`8��"Ѷ	i8�;:�L�*�y�UtGKp������H�џ8�4.�x
+�B�Jo�<Ў��S��b�GK~h>)%�V��o�i���)�گ��"�,�Fғ<�~���hH눭�·$FD���
��QG@�gX��,�a2<����(��R���b�*��"�Fh��:Қi@��	E���ޗn(�K�v�kI�]2a�� @h��xz�EӷYq�������ݔK��.�~Z*���x��iqq��(�F�������d
o��.*Q��8��>�f�� <#���a䉥�֗Vx�LG��L����]����>ǻ�R+��˗�]$.��?�N,Y��r~{�^�5�zi��`\ݐ?k.�p˿!�����o.^v���9�,�^\�7�r��2�C��f���{�"R	�Er�C�^�������'A��9#�Ղ����E�P�d��� �c���5!��rs~���?�<��P	�s�Qj�(��o�g��l�j2�<�q�X�'Q�<�~h4��-_Dx��fad���(��[D5����X_�������}tr�k��Ú��\��0y��k8�S�s�`d�?����P7�Ե�7᪸ \����Q\�*��WPF��S
W�ъ��G%��8նk��o?B/�1�3�����V��_P��a�ek�J�j��j��a�y� �Ϛ�A&=�׏b�l��TJ�
��0�q[�q����-�w4ԯ��J,$ �z������"��c�Va�Dmb�ƾ���*n(�w��!�'�Ќ�z*����%/��2�G&["�;�0 �������G+�
T<�ǢD�_�Z��兠�Y�' �z#C�Aɒ{��i�T�
�
X���T���a F����ź�TWm�DLE0��ɶᇂX�ĉ�L��w�=C���햇�-�?HԔKb���E$�~;��r��i�GAG*��԰S�'��F+���	���q�\�Qa��a��4�2�;٩�d~F����n��/Ka�@rj��/����eX�5��"��y�S	C�N�Y�S��a�����U���F+����Z'�8#Y�cn������?����������Ř������d��R{U`^�{g�%�l\q�fM�7�v��Se�V�R�3d1��}H��
���S��T�$IÀ���<��-ȦG�)&E� �H�Sn=�Է���J�dŹ��8�Q���|���F-L�z��m聉r+&y}~������p�n��iL�@B�S5$g�˳4�����nxS\�_���.�s/�h&Ҝ�Zp��B�e��U�T���VU��`�=H���������g��|88�]w0�Z�����8"���jx�4L	e^Q8#�WɠFI����R�}�wJ���2-����!�.��a��x+o�����oE^ϋ�k\���Pha��*+��Ȇ��7%>E��wZ|`<)�쎮Ϙ��Br~�l���`���4L��+��+�0ɪx�]��#.c�{zZn �����퐃�4S�Q�\���=��U�(��:<:e����y��۠|Ex-�FIy˔K+��H)�t��Pi@�p�_N)�F�ބ��H��`;Q��Y�0*Y��,h���<a���ŕL���5)E�v}E�T�l+^���+�Р�7Tܹe�70�Il�bAĒ�&g}�}�K+j�j��#l,��069b�)*�>}��=����D�Q���u:�7|w��]�.����tk�N��K��hH�����wZy	�Lɶ��P��Vx��\�kڷ�+ɰ)dݧG�U\$-\l��n���$-^��j!�r�5W7�N�g���r'l���鳽���8.��`���\rp;�}�f�#������J.��/Q�����:_��ͻI$f��Y�Tx���*u?zl����f��X�Hd��wٌ��Al�Pr�A~+�ū
����k�}�.
8u
�"X��z�T}KS�^����fF��3|F��ɡ�/���2��p�O�V�`�w~�fK���o9�^���P*�e���|Z�kǅ#x���.ym�0��w� ��U;�0:BL�WӣrYG���w�bHQ�/��+�zNᳺ�
w&��G�	�l
ts�ۀ�����h��0w��$�4�)������VTcKS2[t�����r�>��i���U�i���=�x]�l
�L�殖��<�R���RA��/$�}`��`��uZ �9�"��Y7Ƽ{	�q�2ږM�G�|�!s$5�5�%`4�V05SbqG���l��:p��+�s���+X	��,����ϩ�fz�!�Q�_!g+@�(��J�Dn�w՜$)�j�z�	k�-4�tf�5� z�/ƚdp��t��(�;��HjfI�dx��"ڻ}�s�\�]>ұH˰
J�/V˓�Zt*��{16�i�6z3<����KZGJ����L6� �u`���Xr1���5d=�W�-38�>S�C�Y.�{��Z�`fJ�Wpq˒����A�%�P߷G7��+�{����lS]Ǌ_x�F�8��S=K&Roz������/M��btڸZ��xO�ȉ B�$�Ƕ�Y��S��W8i���`�_%Wmֽ����=Y�p����`���z�M<w��ڵyR�-P~9�*]�Ɉq���~�p�^�E:>�.dpy=¤�BpɊx!+o��6�X� �:���CLr���`��v�'�\��J�<a���B�r��7��F�4��k���=�P�[��8�����U#K�_�o{8$yS`��9�7�&?��֯.ld g�N��7�W�_����1P��]��o��L�#�E�'� ��KaK_G�m��s}U����@�I7:]~0�d[��F����{v(l2aS� ɿ0n�<�`��+��+���SY� �������銛����`�)�/6sS2<���"�27��6$����e���MY��Z$�½��V�b�{+�����@����7����үf۔|��>߸�L��7�"'���mn�f^��؂Ӣ��u[%�D�5E	�o��e�K�Q�p�i%���F��,�*E�oZ��N|&sd�!Mm�Z��z��sKj=�|�uV�NA�ixܴo��{�m��@
)���_��N��4[+ɣ�tΉ��l�mǫ7�����>L*|����ɉs��qy�S��$����B���K"%^�fg��r�X?��[t�H����g Q�}o퇕�j��/@�k��^O}����MтJ�{\�Q�o���50maٲE�������4`�ˍƵ�Ao#����|�>
l*�O�ў��$R�ӱ�Ì�cm��r�r~:���ϰY��Q˪��H�a_�kSX��h	��3;OښK�
�ڜ�����x��e��e�����L�����$Xr�T�Ȳ���	��l�G�^ �.��i�6�}+_j��K����:��g?�[_�g��e{c�9�:w�g�.O�S������o���N������i�_�Ry��<}]K��o5�ݗ���t8��.��g�	?G5v��Mߡ������jm�%n�7�u)��3CE}�a�f@�?ob��ף_�6 5g�]Q��B�O>>�w1S[�y�~���YT|'���V0�i2�����o#����8��vc`/���y��I��ଁ�HiM���>%OT��\b28�KεϦ5g�\�vJ_`�c�N	p�(|�y��&E�����I"jo,Xl�o���;��Y]#��b�����3erB�?3�Eȕ��2�N��;��������Ǳ����+pX)-��8�� }� �O١����Rx�&���W�3r"�������n����R�����m
���H���Q��T�]����>��@��L]�16��`��u����Ӻ���r:��r�<����#BsN���,f�2gwc�����޹�"x�1s��f ��JC����:�x��h�>��I)JJ}��D�v6n��T��;>>G���N7/�v滸o 2��i"~����K�{r7�
7���&������ty��-_�?���K�<�zr��{�}��L{Q3��o�����)E�N$�X�^|�*�t�H��S��u��[��� ���f�:�fb�T]~�i�� ��%��@�� ���V�f���t����08Ŏ�'Oo�?z�q�#pe�@���o����<c���C��%ܨ������u�0dt��R�V�>Nf��c��{/�A<�Pw%��p���2��w�I��?���U�{��D�S�W��T��=��{yg�������O�ڜ�I��z���.�	���������Y��>�^��+�Oy:b���� ���o��'��ss��jQ��#�"�9]o��nv	�F9E~�������^���	0'u��#
�7՚��A�T���/S�)����Dd1/oʁp��{+`�R���;NmkY���&K���T]wX��^4�QD�H�!(H� �h�TA� WiҋR��#(�A�4QP���U"�IH�}3��%��y��Μ���3�;�Ԭ�z`q�Ƿ�d�j�/��b�D]��|���ߠ�9*���rr&�|5�S��Ai��}Eeٮ�4s޴��íQ��ޑr]�"v�x��<�����U���+��g}�*�����uE��/ܾC�������P���<�Չ�09�2~��'fDDGA.�3B�jL%/ ���_�M�v\���C鼖���h�IB�I�x%luwV��e4"km�|ڙ3x�������\�����\k?O$(��#�t^ԭ�h�-��v�7��zo��|c7�A4��X�e<�x�6���A��鍇}��)�[#`)OD�QM���)�^�b��M/�����?�9���-�K1i����Φ$���!h2~�:4F�pw.>N��^X�o ��T�H�dp��(Ĭ���O�8�
�/� ����E�W$������J���bd���A�V�Iԕ� j�����O��+��W�b�����65C}�Цo_�%�u 0;$-y�������۹`KA'�d4X2܀I<G������E�� x���%܁_6�rf-.��;��{~%�~#�P�}�%dZ����Wz�{�����L�9P� 2?ɲpY�,�Y=!��o��:B4���rvMHFE!߸�K�����q�0�K��䉃�}ˮ���@�E�!hO��R�v��B|�İ�j%���ˣ�s�R�&��2��fv�Z���=������"�0K K���)r��0�������McR�&=�����O��)7��!~)>zѲ��xi���d�7%^�J����}=Xw��6��(x���@���r��Jh�ٍ<��rQ�N�(�NA 0□e�Zg�<�|DyS9��+4[o {%Τ�*S�߫΀�n��,�Ҭ���|=� ?�k��y�$��3� �����J�s�)��b�o<��fJ���9����!�
b���^	V���ܮKhڤ��v��Xzg����t�~���gt��rXO�[?�{|Ů�Ó�c��ϯSdM�[pS����֙��z��W	���s���@(�T��ڸ�C۠�	�e�0������D���DW!N�
@P{�E��X]��������,��b������E��_A������	�׳	{� ��Vπ��DJ�66�f���Ok�^��N�zǷ^I��q�y����&�����F+��� ˽�騙�q6�Ͽ�����s�2�&
[%&-ï�.(�����������T8w�zM�d�~�I�A��qưbjV�˶�OS��[/i��*���ɢ�K���Z|%�W0�-�
�/U�b$ҸI�c#2�-薶^���SG��h(-�������pU�h������e��<V�E�<u-���n�P��ҩ�k��haHx�S1D��8�rOǁa�v�<s�C'�>���>_�y!H�DCH@/��؈3�+�z�Տ�(�HuvK�<jT21��J�'X0�ݪ����,5�B���j��PB �(q�;SY%�f�������^���$Q�����ձ���\�)�'���jk(��t��t'l뗠��}vQ6V�zaݚ�C�eg ���P�
�Ż�՟-��n?�]���Yz�j�NT'��<n<��C�e^L$S�_����X$;u��J�ѷ��-��h�n�~���sHaIT�ț�U?�!����`<K�Rr�1�ff\ ��Iߠ#0G�?F���#���>]�;�t��.9����0%7�1���?��"�F��g�����-�n{��tp<�/�0���qm����!�R���rT.K@5�<m� H���+뱃	�9��W�,5?�ZH�$
]�k줷u`���_�W�l�Bse�Ԩ9�+�7Ⱥ�$�>JW�o��_�Ʉo���RwW�+�6wP�'C6���3>���m3���Jw~��������P���ԡ�3i	E/��d���s|6����U�w0g���Y��K�j�˄X̢���(;@r�Z��rWȢ�q6�� V��ʻ\;C�!H]UC�b�GB��ɵz�e��Mg8K�[������0f�s�����H�j��j�!������2�|Syʪ�g�\�Fi���Ct�]��lH-��E�FC����o)N�����Ы�U���ڥ3l3C_�xΕu�-u�}����*\��z�؟����4�v�t�2h($���U�Kg�Fw�Ja��T,v$�����B���6BCw#{���GGk>͆��n6N��Z��^�Q�� Z�6l�Vǐ��_��E�V\�]TQ�ݵ@�^f�C)�[��|E�5F2�-��M��X����y�ڦ:�����=o��C��0	?МJ��A��[�>�[e����#JD���P*S��]��A?��
r�~1�fae�1SR�oY�`t���B����԰�����I}=�ϸI���l��^��=^��.�0dL��ک�؃������N
��/��6�Gw2<��{P�!��ۻ��T&���N_(��s.�@�X���||:��Ma/"�i5���tt�y��JF������Yv�ث~��'�e$b�8NC��Y��z�	k�fS�W�%�d�Z���j�R7`�T�:٬�A�x(%(u*}{Ii��?����V�K�`�K9�@�W	z���1%/�����˩J���U����L
��-�pz��Ko��Y�����_����t+��W`gU �<Bl����̪u�?�'{��J��~� )�%<iV{��rS�L.uKd�<R�iٍPr��a �מJ{�zx��;�=��x��՚{�3��WKXm������R�0\Ѹdӗ���$2��)�o�Q:����C�7�H�@xv��>+3�#pG ���;_
g#g
�a�D�@k\�3��	�ǞI��/��������(���9lzY����Y1� �U����m=c��b��骻����Ep�=)$�:�?#��z'z8�,*�U���v�k(����X����s2�yz��v D���z�*�HK�rN@K��^[��ל��\���Lsb�u�w�)n��g���j���ʖ�Ѣ�*�qȄ��<�,�B�,�b�
5鷚��s�D� �d�j��1L�)�8KΪ(z�=�P>��UX*Lo�$sx�m���)�`�v3%���vY7�*�
c�r��]ggX�~���^�k$�l�{�tY<tI/�2Z�b�=��J�J��r
���~��(��qL�.�7%�o;!�*�v���(��L�OK�����D�h9��{Is"y+�� �H���~`��֣_A��]ٹ�u-*��V�nX���ʼfr�Nݦ�9�5Cr�u]Q�.�S�����Mx�[�Z��$�{-u3����@�bOU��c;ױ�kr�e���@7�����9+s��h����in�y@��L�P��X�F���mY��>h���g��*�Z���<%�Ώs�'άa켖���oJ�Նv ��}��K��r��;b@����2����}�;?g����F��iMݙԖc�����h��"��-N��ڮp�y�X�EI�e�DRR&	E͍͸w�L��������3Հ�=�Pָ��ꁤ����|��ٜa7nΎ�d�E���gI~H�(�����nw2\/(<DR��"tif�wݙq�P�z��GkQ�s�:
�Q�<��;��aeƵ�'q'z�1�E������H�
����,<bN�ː;
A��E�
�˯׵�e�Zv.�(��	H[�z�Թ{
�͡>!`e7L-�����kĐ��}���8P�$�ЊfG4R����~��Kc)غ�R��Ӭcy"�S�bzz��2�Y2\	�:A�s!n(��}�;y
�li���#$=-��6�6w��ؤ�|�W�wxlSmr�Ô[��]3�f_5qr=��g��,��|�l��	dL���L��:�!O��&7,���j�(��(�U�"^��Sz_+��|�p�u�0�;}��M�m>�[tlk��<�6!9>�ʣ����홯�t˓��������P��K�Z;CIj������'��w���\}�T�q�N~���ǳwF4��Pt����L�4mU�i-ď��^�_�Ѝ�zS�C$�����p���0�S7K�&�(/�x�N��l/A3[�_� mh\�-�����h�d�*����;3�& .�hi�	��j?�Y./ŔIr������|ܱ�e�5���_��3�����Q��T�f�eh
J������c7��@��&�HjBdTp��ՊR|�y3�'P�m�L�mO��;q��bn����Y~v��?�bʻ�V��T�w�t+q�lu���Ro���������&�h�z��d�o�iI��e��NS�'�謠�����v~S��m���ٍ���k�6dڡ��̉�H�c�i�ɵ�`�D�2��|���+�#�^�ve�2�M{����� z޶�jT�vY����tV��I�A���@���ho���YW������ �S�g��c/�8�j�5,�O����y�cPv�{���{>i�A��8�=v1�Jถ�80k�uM'ue#d�(87[Q�:힑��]l�������﵌�UY���p�p��]�C��:B���"=ߙV[�>@��Е_FTB	���w�&'Q��,컩��$��u-d��s1���Tu�M ��fW$����~��	jgG&���Qw2о���h����9�[�Z�ֶp��D�X�J*�1(������\�]{2����]eZ˜�{�ɲw��8iCnւGy��[)�ֱ}.�>p
23���-K�����` �=g�_Wn�	=�\(����)�M������w�Y�!�J�FM��/�&�k��N�1�PJm5�>�_{{n`�|N�
�}D�~�G�=mZ	#wP;sF]����ye����pd1j�u�N�5��w���=���6�2��%8�+�����&�8�I�3����!�3��!�x���IK�#.�IE�ڔ��O�?�}��ǩy��xJ�����F8���4��bN�~e�n&;W��Ƈ�o�� 3P�@�x�D�E�h�v�%:}ss�\��>�x�qG|�D�Fy�p� >��M2��c���]��"7��gͼ��Z�J(�a�r��K����w`�"�=Vm���n2M�!��aa��Y~�ѧ�NgM�ou��l�����:�p�$9���/��x��߭�s�M/pn�Z0�(���h�)�_4�`pj5E�R\��������A�Z��3R��k%~Z���m{qjâ�oƗ�LM�_MI�ˢ�\ ��Y��d _�\[Ϛ/�7�H�2|�[�^�������(��l�"��S���X4�,!!�u#�lnvc�znH)�LgzZ�0|�c�xjBM���� yU�מ��͵���vc��cC�4�C�[��/J��;�K�m$���z�ގ40"Ň�����y�;h�*�Rre;��k��%Ud��္����w�H�i3��mEb�|}���eQ��=H}ф7k6|w��W�i{�q�`���Q��p#&m�+�P�U��8�Z����9�J�UM���Z�M��Hv��)����4�c_1qy�=�M���I��nqw����Q��<�$%��q��ʙ���`�gغM����K���R������:��k��-�����qi%��K�W�;���f�w�xX�2 a����c�&눔��5y�,�B%�J�% ��n�CDt����!��O�O]Y�ܘh�c�7����#<�C���+ F��`]��i�Rmjʥ�0�t,����/�-e[�3���$�M��&h�.\�[�}��5o��_�>�$���p���0]\�3󏺱ՊU�6��S^R�ˉ�m�Կ�0���xi�������-F�9��'EJ�.�tI�� ����ulI.fm$_�T}���	�����@{�Xj=�L��j��; ۠K�!t1����� ~�RQ�b19(L�Τ�7'�<~��ĸ����XLE(�v��L�fP�F
�j�۹���#W/���P�A� �0��!��>qS]�gv�hz8�Q'��4NMX���;08Gk�pe~�����iiT\x��UB-}��[t��S2�B¾]�v��}�h�_f�mod�Y��,'JL� ��쳔��OJ
گ�O|��ږ��9�v�֫�y��i�c6I��{f�*�2�y����_3������'��"Õ�[�~����k���7�ӊ6��8H�3s���pé������ծ�s�鍛�)p�D�&��B��c�u��l�)jo_[�-�٨�Am{z���e4Q�$Ƌ�مOI�i�I�~bEߢ��c�[��Ԏ�%$��[�.ʁr��lZ��}ݟ�93F-Ye�Z�h���2Ӎ�1k�З�� \ZZ��/�C�&�i{��_�{���wK�jhSyX��� ͎�66�ʰ\>Y������N)����^TL�k�c��,��p�3^@v�`2ng�_��(��k�� aaHQKlb�J�2�*�6=mb¬��'�	N���򏿳�.^��3U=4�Y��ݱ�D
rc�m�r"7+�*+�vP�ؾ$��g�!��<��t'�c��mg��l7Pn?@�>���O���`rZ �B�&Lz�p�o9h���H0ifm���E�lw�YrKZ��Dŋ]{FԊg�`DϮ���S��tB=:�Wq�%M[j�q���s2���wG#0����\��$�������@��T׈�̆��|�<YP��a�Z�N� �z���r�l+z�,�|VJ��lQiز�~��O��-X���j
�! ��kfS�z��Ļ����<�ׇs�A;��v;[E(Yo����S���-������[)N�d����-�mn�KßoQJTN3d�2�샶K���q]�A%�����w��)���W:ھ�9�E�����3�h�Y�Ran7�������L=�ׄ�[�H�κ��Μ�g6�Tqī�r���K$>k�H�4�3M�j辩�*����>?A������f�W#����z��.������T��0-�B��ƧQ��2_�>�nWۙ��:v�	OOdR�w��6��~�̮�+�ŷ���5�P��~�K���`�7Q��j�ɑ�]w���6&��P��e�ۼ؎Y���-3��|6SR��;�P����'ބ��K9^%M�R�٬��>��؂���}���W(A%l�֜;+�掅k�t�Ǫ�.q��R7�������:�k���]����������t#�"Q�"tׯ�u����d��.O�����P��Z�`�ijP��wβ���m
WV�n�m9`�s�*B��T�\�V�/gsg�o �t�>�슮Ռ�s�H�_�#��N�������'��p�4�~�ěw�����~οʤ���w?���'���:�y�}u�_����O�n��.ި|&��Z!d��n��ʃ��+T�/�d�f\f\<d�>�|�Ju)it��z夾�-�&��SL���w���A;j���A��xv�a�[?�Ө��L��o�]���ڰ3�n$J*�����d��\��@���8q��Yv�oÃ���ݠ�Z�����Q�a)��>���;�T�������%���;��,����5;h�3�$im�U�V�B Gr�֥��H̹�3�������9�%���Le���ߎ���M��|N��:1Y>�y$C[�����o�у�2����$ILWS�����r<g���f��<��%��!ѐ-����$�[Rɸ�+y�����	��ߚ���t�@����w�P:9h
2�D-���`Mi�8	��ƿy�mO�(M���圻�}��/����s�F������D�!ӍM8�Q�d�`��l'���K�2�ވ��/"������UW�试�x
H�~��yg��f��G'�%%��Ng2쯁4����ҹ�9��!�*�#)�6�Q��B�t��_+���ߞLo��*(�B�O0R�au���=qФӺ(X���Ғ܏�蹀/��*����CV�K?��6j�����F���J@eS�=�S4"�%E�l�+5�b��8h��"ٜ��|����]��%��`$�)��6,���b9���;g���f�?�F8|6J��A'�u��#�Gs^*C��7!���a�뒔I�*�ʏ�U^l���n�ǝ0�t�k���UG�����~�ZG�ӆ�Y~]es��uڬ��L1!��PL��wL`��E�YЙ̼O�ב�����������/˳��0K��3%ph�>��,��ǿV�sΙ��A���V��{�A��# @�)�cl>?r�h5N��8Hm��a�ݏ�'@��Q�m�[���]Wy�#`l0��i��4��M��Mq�F 9z�Hj�j�NÈ��7����MN������9v�K�3m���(��Qg��9f�^G�˦�g�i/��I�Si�Q+����_����(.��k�2H�(����D�y����!����k0�tU�w�}���N%�bs4sÊw�d�˖nAb��+t^93� ���
�<f9ױɬSo��*��w����#
C�����9�����\���� _���j��ր�(��>�%%?��āy�dx�r�b5�HI���V�nʇ��߇lp�0�쟣q_���i��f�i ^T�g��ĝe�X�d���`�y隚�9X�	�����{�hi.O������I��cqb��0PA���°@j4Nr	4����ns�R��Nå�?��g�Y�����m�������\�9�m ��{͞2_EnoY��ra6�S�±uq����P�����d_%��,2�F0ϹL:[�&��Cۤ�/Oe�a�:��r�u��#t;��E��ﴁd�Z�uo�����xi�9X���2�W���!��*�UW�S�o5�B��� Ǻ�G����2 Z\�|`9)B��pd���� N~;��A,��_ י�̆��ll��F��r�y�������!�L�|/��&�vQ���8��.����hnT0ޙ�|����4�5���$sr(^�����o�K�U�BH� X�hin�'ꖧ�:��/�r�Iv��A��$l^�=��"Vt�r��SL\Y壥K]�[����O����s Y�I=ۘ~��[��C%��D�'��NTn���A{�	A�B�Fg�Y$�kˤ��|9k2�&�`qn���<�?���V�H'�����/
�s�'Hk�D��t�l¨�N���6�'�E^U������\M���޸�,k�P������BZEy�-�x��3���B��|�����(�t��*7�&p8(�v�hk<QV��?H�"U9O�3�"l�O��͘J.S�^�(R@(���=%[R����IvB���>�e�����˲tr���c�u�|�����=�������= ���~~L	9��l�� �?gn9�~c�h-y����(�g1븟O�6(�\��Cz��s;������ͩ���Ig�j��BP�&FL�O(���͓M�S`P���e��FSTp�o'�Q�/�5�s9���Y�Y&�)�:o,������aA����wQu����Z�{�t�0��j*{�*2�UQ˩l'�r�s(l�#��i�o,;v�^R-���N�H����y��/#����ED��`NC&o�t��K�y"3\{_���z`�`LJ� �����L���q͉�k�c
x0R� o|�,6�SP]�^��娷�Te��zY.@~�;[N�&�n�j{�D
��No�>b<��F���Hq�\�d�Lq�(�#�m�F6Z]�UU��?މ�a�:ߤ>�eA_���+u���?��A����X�8W��$eJ�dE�W,�lb��9�
���{�l��$oh�l.R��O{x���B`!\��f� y���֨����|G�ޞ�u���#���eWF���O�\�t����<]1L�U�(\[��~E�c�ȇ��-c�E�%����e7>�P�}X.�����\��%���s��T)P6M�V�7"2�B����>/�V��5�Z�W����q9<T��(|^�	_�;gj����YH6m �5����Lf9B�B���|�����,�#�<Y�o'��)����D�3�L��i���(�
����<�����}�>����/9�nb���k77h� ���Qr\���R�-N���©FLK�F��W�����e��1�͢���2H@��$3"��L��̣��x"�tY�e=n�U��T�a��
P3Z�?c���v�L�׀�A� ex��>����$�#��uP���e�{L�cCZ_zȍ�4e�=�A뇃���{��ĥ/�ġխ����0��9�a�,A��=�t�3�k�2��Ƭ8-ۯ@�乾ʫ�@���_�Bc,�{���Qwl�-�r���&q�&�u�Ɲ�K0D(���S�
6�����a1�	�Ɲd���U ��p]�X,�+Tl<Q�|0@o��]�g�29-*�9�)����Z�b. ����E�,lT��2$�v���-C^hS���O�L�Vޒ��q��PQ3ڌD��8KŇ� ���	_���A��T�v�,r��ic#z�vȏY�z;�-�K�~?�6X*���%�Na����ߒ��hsU�P�S\��
6���.³H���4�u����yXlzMV�:�	�t("wI�\����.>���Y�C(h��l�ޑ�H�
�(����7��Ӊ"��K���п�أJ�B��t�}��#7�*g�l��!o�z��P�S����xwJ�,��Z%������_sǪ����$�N�h14b�2qV
>��s#�����Q\�v�XpgD��Ж�}e�]��	nЭuL���Ll)��$�������6�����*�����m�e�����=�5cK��X,+��M�%)!�_���k�%45�;4=tl'�R;t�y~/6>Ȃ�����L�n��}��	:��h(z'�V��c�)�����3�!���q�^�#�1k�~ิ�d����bt�W�1���D+����wN_x��-�c:��$�@�Y?����H�1S�2�TKsπĨ	j�\��؏�"$ſu��F�6x`͖� ��[UU�G�����ȵ>��h�OoLqs� �r_��j�����]5(քa�;�$�S�����*��l+g��m�r-���	�fF�f�Zs�ɢ�C��x�f(yLw<|�_�J��G�����_���Ϡ�&�͸#�^Vmʯ�
��:Pw��a�+t���}|4��,��������(@�_Ӥ��lFt��3D�saI ���-d���U���F^~�ːՋ����(Mz�lW��!��0��:���������^���n����O՛��P���'�lp�%���NH�G7|�a��)a� "u)ZKne�]y����	����(qLN�����~6�u�I~Ui�G����PxBq:��d�6ZKE�9r]��d���ha�tv!y7X�`u�Įz�/��#iePR���+��/�ª�3���ud��\�.�i�>Ѓ�C~9�7:|`�	�/��@����;"h�p.gf�[�*q�A>e:�`��ї�5��N�-�_��l�<��Wu�*6�ax�`����c�a;����W�Z���g�6	�>�Ӥp7�d�:���2:G��ot�8�3,nx=�ڀ����@7����Dn9���� n;�	t�
9�w�h�g�T�'��8��x2^�sB��t�)z�Rԥ�?}a}���%(NŇ[�����i��y�T  �.�H	5W%´%��a�z�&��j1ɹ��TNt��}c!�p�.���:Q(S� /�2l�� ﮯ=��ܾ���AL嗶���S��,�0D�a�u�.4[ �N��ܯIQ���P�, �v��Ƅ�Y�����iԃ`v�"������,��Z������`	�p�8ؑ�m���
�I��}�����Z0.�>_-1W�.ۨ�����?�U��0>�N��2/ҝ��`	m���n���2�I�dx���k"�OZ�f�҃< �/,<�}[t��-@)z�e��*p�d���G�Ώ8l�e��z��� u��;_/�Uѣ�5��ew.�ܷmS�W�u�~u�Jp�<Yd������	��+�x����?�Q?F+�}w0yeb�q���s������.��Zp�,�ʖ�]�B��<d҉���=i�f>Z��M�杗1;M)0Fܠ�rr����Ih��+��W���;�0a�@k�s��v�~���(q!{tx��{�_"/�.���<����"Z��W��[z� r��u������⇊��ڒht<?S�����4������������KlE���� oS3#��E��Wâ�k��
@ւ;l7���<	 ^=��UfiFc>#%���э'����R��wu^(ȋ��)�����֗Z4m�JZ]��=�H �қ�>g�� �l�ڞ(���^/������>����N���$�����z����P����u�[����[txc�`�|CSN<�jE�咾���bt��T,Әw�����.��+
�6�G��Oy����?SO��V`�0k����{s	-�u�F�YP�8c�q�4��� WKޚ~llu���eBh�C#�W}�����������/�<���Og��1�U4|�yTel�����v�w�ț})�&�*�ox��@ű'���$ �h1���'=��;���G#���A��?W�t����W��`es��P�T(Ř�wc�$ Đ�`�C��aq����?	��<��U#6O	����z.������Ur�(�<
4�qZ�����@��[�ƥ�z묪q�ړ0@G#�GS�|�cSw�f�]�l���v� ���zP�]��MSSݿ�&��>��N��n����G8Nu�M,�e�Aڱ�N���ew�vpS�[� ��9�?1�她^ǥ�u�X��S�}VFj�	J�������K��s��j�+u?��/=/N��y�싍 �p;��"]��E;��p�dyu6*����QF����~�����bc�/X ���p��K<Â˥��`k"��Oo<�*�3�L)g��!aS�UU��#b�exu��瀨�{A.(�H���ܻ,�� �2����}ێ6�R�	('*��v:����Q,1�79�d�F]�{�= +���`ݯw`Ƨ��{�%�a�8S��
��'��T�gS�@WM��
�œ���.��G�z� �v���t�d������4=���u��,��evڣ�%��"�{ea�jQ���/�]���/��=�4��^��@'�R��2C]��b���6DI����P�~E��1)��r�h��a�*��<A:�[�lD���Zk�s�ౠa��}dk�[���D��	�7�0�����hϭt`72��]M'(�T���i���D�%�;JT�dqOr�Y�[+�	'�r��_��T���>G�(�~��PC���Pu_jG���'�l;��	���4\\%ܰp�]lA*%�n� H� .��B;���4��>x�0$�Z�k�+jKQq��J��������,�M>��tj?��HH�P�}X�ݻAj���&!�~*���P>����E]��{=��ț����s�|;�q����'�͍��Pz�����,�{�y��j���'�P�`�B	~����M*	��M|��x"�`]".n�n��?�H�ã[^r�z�i�~*F�B/U��U�#��h%�
1y�ׄ�T������D �_���Ǿ�0M�ͨ
�ڳ�}�~��-�9/W������^� ����Y����c1�ͫ�0ǣ��& �x�e��g<���Y�U�c���_����7��֝��an�j���ZGQ�����Z�[&��T�lR���f�¦Uk�M9��Ϸ��OR�����(B�Oۃ����7�%��S�7ٛ�jTF'�TSZb��<%��7�y���[i $�@p�5��c��%��n	�VJ^l��`�/��?rs�D�ǴD�I��
��<�r����z�~$����"����x��|Ʒ������-<���ƉP:�=1��^��4IсmU3��wV5;��z|��$�C^MI�D��w�4�yx�$���09H�rs�|ص`��n
��gnF�
o���� �O$�28���!�������3�] ܯ��n.A��2��2ӄj��E8���������V)�c��2T�%� iVM�7dK�kS��I_��,��($&cg?}"�N�CR�G"��?��1�#��~i����k=�m#'���� x~�#�k�H���H)T�� ��b����Ӄ��ā���:�.����@@�8�9�� �~9�B�K�,ov;�k����O�e�b��%�o���|V����@uf����S�s��	c���b�d�a��A߄q}��@F��7!ҷ�}����R_;����[��~P#��}(j���o�>Ãd�eޞ�9V�v�AS�i��#�e�����74�z�N0 :�����V��S(�g{�z�T���PClݼ�M[l�E9�3�X:�?5UX�]���<��I��Jh� �R
�> �s�������SPA�Z�9vͻ?���'�F!��1��A#>O��N����)�M��~X�]��7P1q!�A�,|+���{�fp3��(rU+���4Im�' ${�S�Dǰ�NFS��=u�:s�K�4i>pn�/Υ ��E�.����W�l���)M��@�4u]��y��?ב�Ù?2q������4Y��TU�ܿ���x��,���b
C/��9�\�L��tpx�!�w8�ݑfmo.�g���&���aO� N��y��#5/<�	i�GHڽ0*���q�%�L�	k�����geی�ay�4�T������$[��߾>x����f�2W�MJZ����Y�p���\���R��9lhj^�_b.|��kH�3�vz@k�?�W�Si'S�-������3�A� �8�6L�M�q|���p!�0a�:���h�#FU�00�(;X9>i��o@��V���b�u��Z�!�|$}��#�l�M����vK!'4q�S SX�3��I_��D}
��E�W\�)�n�h����=�\W�.̑�|��/�������:؟i��� /Uד~��z��X=�l�cW���,�ۯ�0|P}���x�sN��`[��ѵ�C�g�]��w�#�W������Ǹ]�8��y����^�:\�Ҙ����F�X��:5'�����z���4W��� � ������/Y���΀?{��Ĩ��4#8XS��_�k���2^}*��?��L/���e&4%�4�mì� g�*�ڃl\��(�^JP/��y���0�� �{���k����U�T��Eg=�6�o�i3k�"T0>��^?��o�?m)Ef�����((U�/L��i�w�(D(zI��7�	)�+���I��� j]�sW�MV������~c���GH+7��2�@S��0U�a����R��C��G��� �mh�{L����P�@n�#%�-i?{�Ԉ׷��H*m�@�������R�7���!>��}�Op����[r�;9���A��[��d�{�v&n�e_Z�A a4�pE߬�C��'��	t�w���Q�j5��ξ� ��x�yՖ��N5ނ9�?����������B�n�+��N��A����z0-��qROQ�5�*�1�?���?���A�7w�t�Jڟ�q��Qh���@�B[$d��7%BkoL�tA��vF긹,:'@9��f�0�3�}R(���,�鯽�ϋ���TV_;~d�q�z��t�$�j=ko.h�X�Dz��!�ɍ�;�/pC�?�l31�Ӂ��9��2�$���\lI+L؝�G5��G���Px5E)�����#���$-�Aj5��H7�����ܱ�Q
L#�k?���[ُￒ4�J�k@��6Ю'���S)��]�B�}@ZMӢC��b˩3�h
)웖}l�{��;5�yv5r��$M
x�~���&%�^00�م ��(�L�R%���xgi�ފ���m��Z̓�;i)'/%��,+�ݨ�)Ы 2�u@��wo�n0�I-�r�Z�� ����f}����~����H�A�ƶ�%��m�*�#���N �>�l�h�Tl�;AQ�B�ms<��r^IL�f���v�8
:�~�ۄ��������z?�`I"��"��M
���X�ݙ��A��2�mbD$T�wTT��3���b��	�fF/	S%���=H=L�7�tK�m4�޹N�(��@$�Ѕ�ſ��*�ȉ���y����v	���Z�_���N��4B�XJ�X��&�hZ۫e�ua9�#2ə����!�%�,����BH�b��ECjGt���|Ճ�)��m27�� �*!AB-��mz���^-��+����7q�C�C���zˁއ6�n�:Ԙ�=8��\+KK�A"u��9�qɚ��q|]n��2�=�`���c��~�MR�m��;�[��|q���,Pv�jN�Dڟ�ԽW�%�p1�cco��D�yev��9~�5�I�B�3Ld�"��}i-���8�y~�s[�|��v	4�<�]m簒���R�A��=7r��eZ��/��F�U V��'ʮ�?���-7�O	+µU�ڞ@a�3�N��llzn~wJ��m��z��-K���BD�w�?w���tr�1u���,R��À���Ԛ��Ȝ>oY����Ly�� ��&n[l�I%sڤ~��+u����o:@�i3�Y��a �.ͬdE��F9��%���^:��]kr;� �V���w��>��=~OC�7%�BG �a7  �gQ����023d\ϑ�[�q����֕{�պ�S^�:EJ6��/�2��sޮP�3~wF��L_�+(�y4S��@b���k�y��0 �\��[���Y��߶0�&�.���A�V�#�O��������� �8��]��v�l�����P�*���6�'R��6�٭�Q�ɴ6�H'�݀�A�����/G\�:���b���!{�u ���o����I!�dm2)���O K��!�*��A׈�CHo�v+)����&�( 
�Ŷ�/h������g/Oj�;�<9�V�,v����@�=�W�� wn��'&�_�.$%�X�K0T��ɿR��M?���WE7r��r��IG� � 1L~� ��M�\PW��r�D�Jf�1P%3Q��5���0M��΄�U��J�a�Ӓ��M`=��қ1v(�кe9�!i�^�J��[oy�&1���騖��߈at%�ϯ�!��c"J�5&�eT�!�������ހdF��p�3��ʪd�lu���<�п8I�q�����f�� �ӃR@'ld�F�^��'���J��y����f5 =������\�_8
���υ�I8�Vs�;v}U�6ټ�J�&�$�q��<�WL�Y�SF�c�o!���I�����J{ӿϕ�^<�@=�}0:�V�>��5fd2\��KC�1&�ˤ�]����I5Q1� %��$�.g/�-dc�E��nl�ar8�+N^?����7Y4"�!PCk�aN���o47�1^l��1�IWy	j(���V�=�@���m�H��{A�@=s ��j޿7���ӳWF��s����Ea=���t|��V�:^*c%�zd|�2K���M���\�U�&�R�����=�t��ÿ ���/��|��j�=!�g�'�\��o���g����f�߹)����j�~��a��85fh,L �-�D�L�F���iY�G�d�B����5�j��Vɤ�H����xř��0�#�[���gؓ_�Q@���$G}����1����=':��<�K����B�GB��5����2��Ltb4�ѣXRB�Ȉ��&���$G�R�4y�A����k��d�%#�gJ(���<)	���qu.�� �%�݂bW�U���䋓�3�Ž��Ѵ��f�}���B:g���ևwO�ݸ�4�5ğ	��Ls	+�����2	��������]���Ӫxr���ga�1r��D�~<��u��$f7�� E�'�������t7����%�Ϟ�$�){�`̡ct�=���>?h�1���?N #�b�� �]{�?��F`JpC=v*��HF�/��O����!eT�ͦ@Сtfh�2@�T��;
�Ӡ��q�T*~��'O����4��X������e��
��H�z��#�d[۾�MD�U c@��G�f�[\����D���C�O�<��8FS�ȂCj")����0ߤ7|ӓ@�x˼#O�6���͘/��k�����싫򋈑U�[b9�O�>�nm�2R��CU�t1am���W3�3��1��f����?��Ɔ�����n%�%@s2�!�!�vQ����2�`����$m��cv�`A��o�������(U�mT<��	�k6ɲ�Cm؋S��L0�4n�*Ɖw�32���Sw�:�s(ö�P�,Ʊ۔�*�CI�wz7eC�p�&�O�b���ݏ �vbg(.G��O�r��G�n�r�-��7]��x��J�q�����V���gGGa��1����%��^�u���y=������$�[t5p����V����/�ѷ�7��0���l<�u@�t���J����J ,rW��w��o��WMn�F�-�}��yaԹD�S6�k�m��0Hlsܞ�#h�(�M�sDW_�݄��`KO�!���"6��n���ytF����f�Ф�����Y�"�KQ��(?k-��kۇܨ�-�,v>�{ `����˶��U��%��>�Z���x{�����u9>r!1xNs�e���ev/��ǽ�^�K�X�C�9��۰��\�?��: ��k/���R"��H.����J��%( %]��"ݢ K�t*�%�,%� �t�7wC�_�s�=�s��wf(��s�7	���'9�vi�X����H�>�^�H������"1q~Y����yj;�|OFC��!H6�;�`�F|��]A��CbDB�Њ�,ӧ>w�Q�Ts�{u��]�ѺS��ܰ4Y�	��=�1��쏔���L�����c�yi��Yw�ƆR�@'���DP���a|i�~�-�i����1���6X�Y��hN�"R.��Nw≡��U$��oP��M��=ڍ]S�v�#n:WD�+EI�b^7t�Qü#	Ult�l��ԑ�F���c!�5mn����5�Ů�{3� J��������:�i�9��8��#�6̈�L�i�����@�>�Eu�}l`���R	���c��J�k!��aR�{� yB;D�7�	;5�sCͥ?0�ۅ�6�bRo�g��vUT��8��ؔ����r�&cI6@�_��O!���D]�f�
U]�(��f&�nSQ&�W-E����.}���c?�f�p��뭭wd�ˠ�]�%��#Ԇ���Z�Zq���~ƙ�E*�H�YЕ����q|L�߼���uJL��h��PxVK��v8��n�eu�1��:OqI�����a8����lG�i��Q�交5��\N�g6�~B�U,��C����Ǹ�!{�w�=2_��	n!�'sd�T�x��Cp$�*�*q$c�v����qj�� �^H@_mmKt�Z+�|փG~Ş�J��P#�?��qj\F ��̫�O vf�������F�����o��8�0���I ݰQp� D3�=I�W��z#@/ �_��C%��,Ф9\�&m�ՠ�	,�'k�W'�b~�}Pu�<�;0ʔ/���s�D ���t'�u)� =
�Ylm�pd��HB����N〛�W�������Uj�u�y�%����W�X���<&ۥ�VӲ]�;�+�&�Ʉ<�5�L'3g��l��B�Өmr�z&� ��CYmM	��z+�ۛH�yJ�+�����F�x}�J�l�����*w������x��ä������m9T��zik7��ÏA�r��_*A�i^ʪ4o��!�*"O� ֦��x�����1�� �rq3���cs�{r��(�Rq0�P�nlc���wb[�m����D��ʢ����mV�MSl�.�Y�Ì��=���o�ѪK�12���8�k� Z1�fT�|�QD:�m���;����"H6�[�g����`�Q��C��;b�������'�..���� �``��Dx�4�"�H�B�Խ7>ON���7B0vX�ۆ��� }0�Q�zB�ּӮ o[��2�j���)�Ü��q�W�G*��v0@km�MA�שּׁ(~d!�����{R�GI{��8�x�Iu���Z�Y� o6��d�w$�7I�3����/�ɌvMO��?�j�'��a��)�܌��['D�g@$�C��{�8�(��e�-�ݴ����~}Q�� }h����7D��еH"/S-%+$�t��ZL��ag?��p��X|���(k����U-��n5<�񿕌`�a�����RZ��(&�w@��n�ŕ����9P��:p��+9=r��L5K>c�bP���܀բ&/���NO���D\��ӎ��T�P���@�\��˱��I��u.#<[�vu�aܸY ���8!�7��;Z����`���jT�3��b?l]��酏-�������Pf� ��1�^C���c��l3D��2��Ԉ�c��c��f���?<�҉WRs�
�3�w�Cϭl������L',��ޓ�$�p�g�<jl�н��Yr�h�tk��W��RȍIz%���}1a;�?�M�񕥷�����"Nf�&�j�r���%����RWX��3if#�0��mr�?�|F�˥NIdo�μ�X]�u����Ҩڭ��V�f��ٜ��wh�N�1�[uӂ�Y���rE>��K!�2G�Gn��y�Z�]�BN���Fg�;�iEO܌�l��%�*��B�k��LFH���s�`��\�����Nm�ۚ����ZLh��(��'R�bKH�[C)ŭ��]�1hA��JE��6l��%���6�~���f&��dG�.�-���ծt�SO2Xte�$�Ͼ��������pnZwj��,3��e�rKwƻX���PFС����PG3���v(č��?A�k_��5�Ԭ+vtw���7$b}�WuD�}��$�@e�e�ᴔ�:`�bg𴔣X4���MEs�����tQ��>bzz�h&-��V>�@Z/Cd�!~���Z�(:��?�`,��fe�Ed��\=-��z�����l�~�;3:��W�Y�'��>p@92��z��w�Թ�ƚ� j�c�.��i,�`\���(�>�c��J���jT�
8�y �M}��2C�#��9O<C����׮�V��7d�ȡ�T�E[u�9F��ͪ�^���̚�cNL��{<o�$,/Zل��_�-Z>eƻ�J�v���K�m����v'jm$gznѪ�ad��.������뙘bg� Q���>7��gE�E�X���d��k`��ȪC�����YA�Ze-�Et���^?�����w߾��;"�G:�eH�^}�WC��T��3�Lw.t�����JX�w������)�k��F��H��������59�g��~g����T��j-��l~����V��s	~�SK0��9�SɎ�9v��~�G�-ۤ�3��������p��S���|c��$?kRS� FK�.����3�c:���)%Cg��!�ׂn�/C���������T��g�km�u?\�֝�~⸳7u�J��^J�����f��@u�xT�N�����JG�!(�_պ#��NZ��L{I��x�9�#g1�9�!�!��/���\#ߣ�L�:Y!c��F�>r�������=��2Ci-e6&J�$$o�B�l�_8 � ��B�r��?�Y#G��^�|��?��d�i��HIIq��J\�OR�v�<o��U�B���M����&�����%�\Ǜ,�M�B5��+�?v��}���� � UD,�"熜Q�P_��;u�Mգp��X���֐�^��7���R���VMs(��������2!��Uƹ������)<V��y5O]fEr��\�G	���_���Opp����O�f�3?��_+����.-�t�q]��>���`���t���k{{�#�E�d�]U-X��8�b���� ����?H� Z�b5���mJݐ��Rtߤ~��Ӎ�0����.f֧�93�'�	9O�(P]��ΫW��H���(���C��*���y���_U8��#�p�&�ApP{Ng]�`�FpYP���R��v�¹���"yɖ:*<�D�G�ѯ:���4�f��.��:�֝�W�AWz�ZZ�kj�Dɳ�<fh�,EFqX<��Mq<�N �������;�w `Y{�̅b=3��r�]#�%���lh�q	S0�H�.���N�P1�0��,p� �޳o�n��!1��-"�@X P'����!��ZY�Y2+�[�c��CXP�:4�oo�Կ����V{�<�Ŋ��xH�?��ݱ�[6zB:����"qL��r؇�u���W~x�:��T{�9�i����~����>ڷ�����\6���n��dV19��ܝ�\�i�}*H�w��@��cr�2�_\�=;s���<17Mi�O��AH'#��p�rJ���V���1�g"�E�gk�O@�jəו%�����A����<�`�*?:��y�_\���Ä�e���4��}��
�@ꗸ�Y�)(�|���R<;k�F�:�\{�;�ѷ�&ڑ�H�����&�/�<a<��fq��ZD��?m�2�R`S�gR묁DJm�����4�-�S�f�˪2-�
ģ�c�k���	�ڲ�N|m�%-(/s���#��t��A���u�n{�|�̬�}��)*r��x9#��}�2~���������Q�(E�m\��	�[���
����]^�rr�[��g��HgrhǏX�Z�-��������:7+D�G���.;H�%����i�0X���]��eof;�Z��G1���	���;�$v#�6�<�ר�1O���h�)R���j۩:�{�]:��2�f{�.�Be�	w�Q�jE	2RE���|�L����tI~��)PH~�C���Fr�k��C�wF��Q3�rɔ">t8�s6:l��S#<m�>�s`:X�g���z<s!G�~��>ԞƸ����>b��%-ܦ�"�#F6\M����Q�xNK���'���3b�^ِ�4O+���L�S)uR��{�f��߾����2*����n+!x7k 2��XfT� %B�ֻEGǜ2��?BM3D����su_���+3kE5)>�"�>�^�jQo䇯"�2��j��J����ME�]fa)��OL�$=%@i���O܀[�n�US�<(�O����ss���P�ʑ䈭@���d�k�s!�z6�T��rt@�N]�xAK�Z�?%o�8��P.t���8��.�Ãbm�E99�	%�։Ěҧ ~�f��� ��z��>��fg]��ڊ�����6�&M����-b�w���Ϛ�ৗ�ܰ<��Pe8̰Нuu��_�l=�0@�X�zQ���?�_U�������xV˔Z_�ԷZ���|����bh��
�u/;=�1��1i�d�oEG�Gq��وDP��1�s�*�A��b4 �[O��KC�bU@��C�r���J�����,=3.*C�;ѩ�F?�YV=������b4> �d�+�l<�8W=��&)��L��T��m��_���Ǧ�tl���3M��Ʈ�4���r���N�Z�6U`����TkscQHH�M���J/�j�'�C�Gs�|����9tς8/h�Xl�8-n��^�HA$J;�B�.so7�&p��"\���S?5�R��Yk�n�
�Y��TF�S�%����9Q3�t����>O��I�}��z8~�PG�u�O�4��x}O�&���?��$�Ԗ�+�Sw��\
�I��#�E^*'�u?�*��'#S����[�#��I�^x��1��]Z�o���g���5��~! `$���Y��a�X���F����Os'����^0s/I޴ALʼX`^�r�7��~����C�'q ��������C�hf�
K��B�Y���WkiZ�Qkk�Em��̩F�Wmb���g�	�ϣF[��,u8*�r�y��W�Kf�)<���lX��뵗����.Q4v��$~lƐ���<+ �kjT��b_\*�ï�F��%4��^<,���ri��Wޤ`�!���CYH��m��T
}�(���(�x[���,�-y0ax��ޮ�<Uh�H�pͳ�#��5��8YQ�H�=�8�r
�Ui���NВ�V�+��vCed����:�MhdE����b&ך��c=ru��S��������f��	"-Z��cB�ң���s+:��_�4d�t��'����"(_��*���c)4kя��m{h*�_���3]ݍW	�
4�7h¦hK	Oe�\j�V����D����e2�PJ�ʐ��b��TV�/�R�,�TS�+�]�ӑ�ם�D9ԧ
���)�Oň'⢪	���C�6�/��ɓ^]�Ma�.7d�6��۵����m��m�����O��d��TR���� 8��o԰r��k|�l��`�)��T�a��d��&%�G�%ȉd���u.M��gx�������ԏ�W���v����q���ü��$ �Z=�0�D�����[cx�\��y���U��h~5�?@��c�Ȋ�Fw��{��Us��g�X��s�w�i?u��/�q�-�%H~����پÃ8%��J��佟��V����	�>��:����`�M�N%���S�'��@��#��_>��o��X�}�X�n�&LRpK�B�ǯ
�(3���x�وje���z?�Ң��<{�g��z㙆\��������0H���w��^S��Ϫ<������e� .�����.f*R	���Y4�������c�;?Ғ
� �H�➨"��4�w1��
����3��Jghڗ�R�K��f�P��|��K`usF�υʭ��1�}Ø�����p��Z�<AD�Ǖ�Pp��a��Ԭ�V ��p�O�1p����|xv�:�V��c��4ØP���\i� z�������?@�ވݤ.ɶ;�n��V�g�<v�Kެx�i%,�9���M��z�Ӟ�m� ���b�8����qK�`H����O��[,��&�r����+g�Bk)|L2��A�� ��-�Bh��u��\��2?
L����B\�w3�z�/ +Ɵ�L7�f���g�Z���n����i��C_�ߩz�
n_ˤ}E�i����(
�~����:w��1���u����"��s��,�W��VA��@���	�z"HV:�a��Ɵ�vg�j �i��y��}�ZY��Ӏ[� �ǹ�H�ܐ���o׉'���To|U�?*}A<�҄2���1+U��⺮�N+���-|p�UEJc��$!w�yx_(a>�'��4-�+AMMl�t�'
j͢�|a4��jW�u�Mh�_`V�D6�gm.��!(�Z�̀���G�3�T+A��+닽�J9�ի��V<�'l�aB̀(R���	M�M��eW��A:����*�,��.%�ǂ:@�]P����t1^#E&t� uâ������f�\��M16׃3���'�:[��� �O��_B�5�)�����'i�CZ. ˿�cR��u=��p�-��^�
���Y) JG3��CQ�b�6�'�&+`�8b�*:e�ں����3��Ccm�s�.���A�E�(��@�p��糫���L��{�LHj��IZ��ι1�2g}'/�Ms�x�q�n����˲�<�8e�YW.��`�SQ�ȱ�&Kf�ĉ�ؼ_h��/_:�����[�Dm㒄����⃺ľ0�=���[��p^x�> �=:�j#-�1���H�j�oBG��/��� �	�M5	��6Uk���z_�����H�
�GT[!&Y����OŋM�s����1�Ĳ�}�Dj%CF���[~H<�y�U��>��T ��N�M�n�'�w50�a'���b���8��.Y��f$9�(N�F?�6��j
�6��ػ/|��5�����B����:i���|J�+�{؞�f� 3�G�RZ
�SW�tT�:vsC`�s�g��
�h�p��a�`sLa0k2b�uzP��N֝b���)`lg�zcQ�E�Z_��?S��
���M|���	�Ӱ�ee�����)zx�W�
T{o���E��W�.��v�>{2��ds�WA�_>�����k#}0�癣�Ԅ]s'K�c�s?��m!=��'��N<ާ�Q�����IEB��/�HV&ƦH���d���Rjx��-ýg�}D��������8�]9�)��u`w6MX1��j9M:��h�8I���qh��?\��r����Y+&n
�J~T��h���7J���~C#&LX�AB��\g�TTY�-��:XF9�j���.{h4�}E����ô e1�=�ύp**Y��ǵ���cH�J4.�0��c/�Y�mt]SK!ř�]]�0}�r;$k5gO9�o�Է/����e�@~t�Jݩ��F��mZ���z[?��j.��?)R+��}|�����q܇�$��k��_q"����@h�ҤU��-��4�ȯ�2(ZՔr/ߛB�=�^�SYE-�iR}C|U��=V�Ch��*��q\]�R�t(,T���5v͓�,?�e\��/��1���}wӝ��ƫ{)�)���Fd}22�^���|����bȔ+,��k�
��s�g�X~(ǵ<j�.z2�,�aEm�~��L?I��]3Ex��;����Ͼ;��!NL6��m�^37)7�	���������{ݴ��Jd����k6���^��%h�g��d��$��զ�W�����PF���/�R1Ec�t�#��73�qZi*4S1.��,��t�̝:\���� 4	FE"5�O��U�PD�oϋ�v�e5�À�5#�=�8u~q^n)E�il�W�d�Z��os�O.�U�c
�Ԥ2���[��"3$@��Jz#�A�s����o���WSnirArg�{�ʌK?��{Խ�����Tw�RX�p5?�ų�����&��Jf��K�{7l�%ngzy���c���3�ã�_�~?\�R��r���@��[=�[ ����n����@h.K����MѦ��Bsޮ������� ���;0Q�J��0-�,Յ�N�u���l� W�Ҧ�U��߬�1�*���i�W'�JM_�k�� {O��S�n��n
)���Ǆ�{�c�#b�ߎ�d)��>K-���J�U���p
Q�m.��gn����<��`c�$�2�"իn��,3�m,���d/�����^��JC}�Po�$摫P��0�ݮwkԠ��+c�?4����(�`*�D��޶zGA���T}�ȹ��7���-,r������!�z���ev�?��_�tCfʱ�{#����)�\�ʚ"��|4�d�A
<�stp�V�,3���עc��w��/`��
��,04Te�Ua��t8��奜j(�^�!>����SyP����<�j�w����p�u�=�q07~�;󓅣Ħ��ir{��c�Yk	@�|,�1���fUu�C�7i
���L��
�H�h�-��xdi��Z��
$�wW��S
�/9���Zw!��QJ�Xf�=�y�8mzA�}�F|VA`��~
�YНȮ`�O���G���(Q5��e���-k~�9�,����V�;Su��3J����3k�O籬6�\������������'|u����i�{؊¿�G~ &�X��;�r��`#9�����~���h����P���	�m�*�����8vs +���PMP~b�Yћ#�e��m�֣�����)Bw1 mgֲϯ\ L\?k�s^��݋Q�K�K��/��Y�ch�)x���~Z
nz���6��Tv+q�8;�B4�s�&P��/P���a�&����A0*
]���O��=$9[d�� )y]��$��^ib��g�YXU�㹝��[�y��m=w���\x�
��Qiu*3�,�%0�iu�{����E���z�g[?-Ƌ��e��{3|AzKK��j��u�%�w�5U�q�R' {��IXg��
�1�!Р|?1���r#���EE�qɭXS3�q�(�{��V�'��PoY�<�w���-A�p�A O�%��c�Ե�F_1��Ef�����[�Jg;$z�
�������Ӕ��m^ p�NSȠ>�Re�[�Hd�?_BLov'�s�ep�+�*�y������ƾ%��d����w�!4�gZCÈfw�Y
�Qi�}�F�A�d����i5F��0�PW�BN-hI�W�~�H��qm����x�Lva�tK�:kq6�@�H;����K��b�u��O����v��t��(K!�L"��t��6"�6�x�L�'���Z�ev56f�?Öc�L��)iZ��t������pFX��3[oD�N��s���~}!�E���ԍ�uq2[�6��o��(�$�� ��_���f��<��C�M�4j���P�ы���7�;�%���ｅ����r]5S�|�pI|�)�@�����_vՈ})V��_��^���xr5�S�<��uM�Bu����X�}!���;KE�:����ӧ��L?0�m4'#����"6��`p��7bFR���3�//ʔ�z���Re$ߓBH��U���40'�	ӔN��o������?������C+�ϥ����a�Rot�����s��{�����=���� 5�?D�B"�L5a��w�zocP�w�"�Ŗӛ\nV���79n�t/�u����S�RRқ��Tz9�����%�溬>J�i���;�R�cMN3�\ci^Y8~����F�L��}�X�Y�Ŋ�F���h^(M�?UJ<'��#�Ǹ�zmE�>A<����9G���B�N)J�L�v]�Z� F�-='�$�T��#�ǁ +t��h�����'�'������d��˲�{�ל�t�g�n��ޡ,�"����؇Ky����d��@���H����gU�5�����:���Co��1Y+���h�G1 F}3�KOQ�O�D��;�@k'y��0��7�#��^��~��%ibW���&t��3�x�J��	A˪z�oKwa���@��5*Z��,�c����No)6K(U/8�6Z��#FAô�I�$�Eh�_���M�~<3�G�0e^�{�3�)�;��R��G(%V~�i������*+W4�`%���Su))�� OH`��&v��d��E��U\6�}�Q�+���q��.����{�<��3�YD��%JR�Դ��ɱU6���4�c;lY�� W��Et�Z3��3���9S�Rg�'�:�Xd�e���zt�%�m�Q����DJ5*��������jc�bfs��<l�G�~�H bI�ʣ
�蒹s� |i�Gɚ��l��n�2��T���at��p)Z�9�:�.��z����4�<�3�b�n�����Ӷ-ýV<��|>;�w������X�����,��Y"7f*Rv�F(���FrV([Ϥp7V�Z&��㽩yj��'�Rɛ�ب5:�]��5k���	HR���e|@9|ߠtv��i!/�Z��0�Eq�^�8�m`ے+Hh\�*[3 �d��#��_�΄o#��߄�4t��nYOl	���%��o�f3~$5l�T�W��1�$�LĘ
!=@�D�'��D�ޠ����,�W��9��\�ߙ㹵u�ǰm��^^�)s�hcW�����P�a�h�纒:����̤x�{O=����gj��������D��xq���F�~kWR�J7J�9q��jm���;�Z�펯����W�6�S�^�[����2�������1BpM��A{S�����E�b4�H���t���8��'u�p�D`\e@d�!�z��a��|����d;�Y��]�Z�ץ.m,!>,9X�eS� �s�`:W{y�n@�!�b�ö,b����P�� 	8W�����C+Y����w�b儞�-K�y^���9������3�?�WN��TB�4���M:ԥj�AOu�YS�Qt&�#�Ѝ�^2]�����:��5m�]oa�zH#5�]���T �M~�xm����!�9�^���JXА8ԟ'����P| [%��!D�}=3�c�P��+ 6֋U���Q�G�(QǸ����p����?�SR�xybq`�#0f�z�z�8p�{$�o�:�����abJ��k��:���s�ˏ��"#�Q.�X5[�w�j����:�{�¯:) i�'�w4:�7��J�����_O�,�8���ϐx�p�+sw�t �;g���K�j��d��w)Sڳ���Q�Mɲ.fS��d�n���]�'xW͙l!�!˭s�^�be���C���F� ��)1��z�t��
*���w�xd��>��2�`����Q�[�����e�B�ٚ��2��R���L��z�N���,�?��m	�xn'��Y���<a�yެ���M&%G�<J�fX�s�9���-��������d��FVP�#�w`�]�8���D�@�(�hsx���F��#�����T���W���#Y�#���j��݀��;��نV�#��/�/~|����U�x��I����k�Z��;SL{��&̸1�T����C���k�kW�n��wĊ���;KP���N�N�Ϭz��P������1�c�U�f���e�C�*�a�N�Ä��{��M�lŏӆ��U
b�9�uT�;���*j�m��5���tğj�>�����do�[g:풚�Y�����8���p?<y�M���V�	Q�)�:e�U�o����~�>��e�=�5����� k�&� �$��)Ƀع�h�=�n� KN[>�t�����N�]�g7U��n�1br��gӠ�b�:�7�5)ۏ=�Z��)iW�o��^��x�"��Y���#7�;�LLtG"0�#�!�|��K!t�=^������U�o�5?hf�5�?�)���sJ�K秬QsNG:�[�0�l�(����֤����f�4׽����&t ��KmԺ���i�f-��N���G��RmY��?>`�og=}�?��f�Ӭm;��k�wm���!����{Kf2�'F�tF ��[{�j��r�|F!�W��İ��}���W����Ab��G��_��)�gq2yJ�a���hF[+`5��"��d���7ͳ9����1���8��-<>1�<R����EQ�>�,�����&L�u�ެU?,h�t� _ưI��\���l�uG]�w�?�2���m��y�b?f'-�;�&�Y��S���H���u-S��ͯ�������
��������ؒƶ���&]�($��n�~;���q�/����p��<�����'�2���|Z_�͟�0ףJ�{5��@{;�iK0��LF�-��qe�C�	��X�kΕ�U�`~�p�~�K#=�,����̫Sr�'jCJ��Ŝ"�8J�c�!p�'��w�����V%Rt��T��s�X�bTc;�N>k=�Β邉�ϯ��Ŭ�..0��c�%�)��s	�_�V�å��7Ƣ����~�Ӱ�\Px@�t�Q������+߲u�a^�N%=�dՠc7bnB���(?A�z��	�'']q-6��ϡ>)���'����N�*c|�z3J8:d�ޏ`~$!h��w����6V�J�\y�
,�i�`��a	�������h���؉��
,J�c�蜊-9�.{�I(�߱��ȐH=�ё�gx�|#�{H{�a����s9<��"���*���ɰV�SǼ3�g6��ΰ�/�w:0��.돴m^���7��<2�doG�p�'e��G#�;￪���t���0��K�Nd����w{]�B��|��F�wKD�.p��Y酵tX5u*�k5���R�n�]?d���r�E�Ku"��@�`FM�I�ꢸ#����p.aN�3��N���������᬴7Gƃ7Z{t��F�t%-I��q�X�6?@�Jn�yR��@p�@�OƙX����L�ܜ���1���K��G�Vt_�P�N��Ai�V��;��:��v��ۨ�7`�~p۔L���	���S-<�-*��#�2��-�aC�4��`�t)S��?�S���O�N��`MG�����|�zL=��'��40ZY0�z�F����0�ɧ��h�j7y���Z`r����VŻ�2|�%�D\C��<s��i(��U�eVV�L�׌���軓0y�åWu�Mz�ޔ���<������D'��Z�@Bk�Ƨ�<F1�`��;-�[i���A��v��֋AB@-�s}+=�,��W����#�����l���5���3'��ۋ��k����Z1g����R����fO#7� Y��!^���צ���<�W'w����>�x��W[�4cVz��2'����8�����z�3�b��J���;���3��n]3ջM��Y�{�x�t��w׹�W�3��#��t^WL{4�j�L��U1�)���/o��o�j��}^���å������e���`6-��ݵq7�DGv�;*uG�(x�'�NΗ3%y�e{�)���� ��H��(�O�ޠ�:��t�[�7�c|�@j]X+����X��3z���M�����L{AYs�� ���5Ͳވ�9�I�w|)�Q�pt�e�5�#,��S�"�����e%��!�'�aϪ���6�+�:�e��ȹBB˽��gt.+�q!9�B�q��4������ ~��>���2��	t��u����v�zQ%i�m�4ji$7~�9=���5cHNG|5]��n��i8ظ�~��Fܶu���L������paİV� ��g݃KJ��?L����w��O���Ӊ��m{�T�Dyh�J��&�6�x�6�L�-���$�����j)�h��ԚY�v���1�p=��~flIF����0~�)����,�!� ���w��LB'i�e+WW�)x��#o�N�MR���\��ˮ(�,�jם2ƺaԸ���+W<㸘ܼE6�l��n(���/-B�Y_y��m��H�Me�`�B�P� �|DCdj��_oj�F�y�_�?ڭ�=\��^6ɹ�V��ps��ߙ��G�7ĕ[ji+%��F�m/�.�Ǚ��A�I�������w�>j"_6�y��|Co�4����ޡSNi�l��u��ɑ�Vd<^��Չ}�7�B�Q׻�t��閨�{�k����'�Gbj�3�U�z��@�^%A���ʹ��=�o���T��u��|��&"^B�D9�r�G`��׶���ȍE&��M�Z�����y�fC
�G�����������GY�x�/����/�|>�"��8�����ۧ4��h������UW`h,��~�kHT�����E?n����@"R��;���F�����#���;8l���9(���E��c:��,ϯA�H���7?΄�s��ik��:�	b�T�?�:+���X#�O�h?�#��S�?(��S]lR��#��U
l)���t_F�8;��-����V\퓉cVA'�3nx�2�YڻU$RN�.�y���1�w�����o�s^<�q�h����7\N�a>T�2���g@��_\��D{��pl�J���ی��2Dc�^����h����d&�.95�-��\&�nBPƗk��l9�#�8�{\�a9�P"M�*��rh;'���F�[?%���{n?4�����O�8:�S�cM.s�f:j2P�ɍ�`��XX#������_i�����IC
Hi���iRW������pD�kd�qr����<��b���uʯ}��^�p��#m�l��3+?��Z�uY��a4;�� �>/�y�Kl����9u���H�Q��\r��8��}������_�C����f�:9�jJdE�S����v}{-/�+\}�^� ����\3k�8�x�L(F�~���8�F�8�}=1��)�����.�^O,�{S�:>�t�D9�l'ᙀ*�_9m�m��'�ue�Y3Jl��/�R��*�N�$l��å��!�,�*���c�
�%R��F��a�娾!E}C�7���-C6K+_Q	�me9L@��޽��1�y��0-f-?�����h�;��I���X��(w�/�N���[�w�V鍭XD���@3�l��D�c�)ok^̓ZZ+�R�o,�1�j�3M�-[;B:��4���Ү������s]ҷ �g�UT��
�Ź�����c����E����2z�~��K���Rk����|Oc*Чsi��B�,��4���ucM,��$��d@:{h���R��<dF��M���ڍ.��ϟ���ĊC倕X�nӿ��W	��,�^3}ű���@T:ڦ��-��y(J�f��(��r�o��Ϛ]��h�̧�*�5���S���W=��&¬�!z��n6�b��l�Z�hA��%
����kZ�����Ȕ��򯇆�����Bvڽ��6���A�3��l��33��*0�]����1�=��+�<����]/�k7ǩ�`��jq?L=��N
{�hJ̈́i��	Z94hÛ�Ie_&�bj�S������o^������>7<��@�\�B|���Rn;�Y&�eꎖ�B�l�����C٦�����g��ó�QE찅qҹI���\%�=E�PZ1M�6F�m�I�ei���膩pȅ���JH&��LY��yQ���D�E�t���n�	�K���X���%��3�<��
k��Ty����Z�%������ ie��>�}����0Ϙk�/|'z�;� (��rs���kx��;`�&��~R^�~j�'���Cd���K՝�����	G��_�h]�P{1�j�`EI�n��8,a�v3e�,��������-�
`}��%�	��]�F��L���!���(����hQ�џ��-�7S���b��Z�:�P�ǐث�t0:шa5<@�Ga㳦L�b�GgX5Kܿ�����ҩ ��bڗ[7N4 �����!w��U�l�ó�Ӊ@j��a�go�,ָ�t��W\�������8pz����wlC��F��l.ʅ���(���������0F��b~�3(n�N����w��5�.�O��Z�:ъ�A��-+NaS�����Oa\|}�锪�1�����(��g���h���8�D׬z֛$�F�?\�G&��k����l���\	9���5��%�J�{�}��n�`b 01�I�]���I��}��Ro�p)W�ʩ�� ў�L�mˉ%���'Uρ����n��jʉ���fs�L�)��Ys) �}d��`���Ֆ����p��7`���ӱ��Os[�Ŀ�?T�19s@l�+�9x��m�j�ԭp/I�W�
'̜II�g��1n]��l'�&?�;�΍��>T�@B.���)�3�x�7�c#�W�G��ƴ
W_ǧt'#���]�Qɔ����A+۱ڢ�9�S�ݫ9���U^qޒ�ڨW�*�ok���ҧ{s<�����ƭѭ������}f%3R�6�Z��8��ɭh�`41�ga���{�}�۫��׶
n0�q=�>�WS��m����<��t�~+���H��r\g=M F3�<;�����S{��*���h���,j}-��X�G��NPg+����	 �?Wry��X�4V�{'N�>��8�o�@�����9u���L0[�mkٌhQT;�"�Ct�QAi�9(�--�-����.�Vݨ�j2��(���MR�G�{�9m�"�II����������-�8�V�M�$j:˥���@!;�9p�М��k�(��w����-����
�a@&�Y����X�j7���<��H��,>c��������W2#U���-n+���ְ�;pV�)�AT�2
=���*(��x��?���ֻ��O��;Mາ�#> �J.r����7������^U�;Ԭ���BKIR�r��)��(	2�&{��Z���ל�J�M�k�7���i���C�)�K|t��I��/G91�X[GF*���7ڒ�1�M��H�@s�# �؀�{�|8������֫�[��ڥ�����3Z%o��ӧ������ǅ��w��ڏ7�{���e�#�YCV���'ʎ?��y$�h�����R8⁹�WpT�OSe]h��S�D��csx	u�gն��HE�Y�F]P��@H����Q��9pSd<��^�7�^�u
OUX���G�*+��N�����Q�No~:{�u��	-+����C�F��X5�e�,�P:$T�M�f�mh[$�{����
�~���X�;�=U�%�~}nj0b��X�>���[�4W�JUt���	��+�a�Vv%M+vת�D���[))53zYv�9�֨ �ݟg:lB�#�?9{�����S���K5=���뵊W��⡉����i��i�p���q���h�U-�{6�_����k��Wz�V��yZc��	�L����3�`l?|����ܤ��;�1v��鑝�u.ۚ�����\��B���a@V1��x	!�*F�L^4�A������Y�g�=)=�YJ �˗W}+�=�Zc����MmTC|3���G�NGjw�[5��M�b2�#��]�d�0��
���/�ߞ\p��>��[�%�w?�@�5xk~��U͕��l�g�b'���1��TQ�/X���V��&�E��9���U�ou��z�>�$�m���=���7��wm����t3�=�F.+ߎ��^��-�]�Qs�����'RxdJD �����9r|�쩡:�}�]!���a�lN(�!~$Vc�WR��ࡥQ��h�p�.� :��} t �!8]��[8hYɢ�#q��<���)���=�:/�`2���lʡ����lzм3P�Cx6V�� ����*��uK'���dU�6���iL]�T㑹hے�ے���?��;��=�7�E��`��HQz��RU�I7R�ҥwB�*��"5�&E"��@(�R�& ]J���&���w�=�q�';;3�2�]wY����b����p��������ikHh����Ms_Z�dxz٠+��A��@	��E%Z4	���V���ރ�7o�-��T7�d�o�ε���1ߞ��`�~� ��X��u`��(@@��@F�^r��^q8�(=5��n��E�hŬ���jbp�,K������Ί�ڔ�x�Lّy��$I���.�O?#WreV>�S����^�e�_P,Ӧ��ybn�1����9�X=Z�`S��^xv�N��dOq~�i�J�������D��:��E���;��	"fq�%_iR�X&T���Z��[�k�������DΩus�h�T-)(2�v'�L?lS1(<�/�^�y{���T��m�L?���e��>�)Q�w��Tc�I�"���o�Ϗ�X�&Z:S��-�d�,�&�.�����i��Sڠh�8c9�����@�j���,n�&����Y��F�_�E&��?^J;���}�aܩ0`0�����F �{(0(�D�ޘ���3iO	-c�OSS7���q��7���EMXA�)��FJ�ݨ�Z4�T��r³��Kk�mͣ���0�c��g�k��l��P��U[�	���?�"\H���Lp��|����o[��9���P����#��H��a��s}���m���F3V��<aۣ�2\��(Lz�+\?l�� ֚;w6��� Q�?o�S0�pF��J��k\�Yf�K~��T-�ջ���1û]�_���6ߛ��<���:Z�o��������j���N����z�������d��n�J���B[�(��_(��hI��A��z
��6>�8�)��6�2)R��(��e��Z�=���1f���Ğ�l_)���Y�1����v����M�8�����t�n�J��3�`�2��-]�Rж��U&Ƞ�5�yG9��v畝^GW�[�*�f^��������?����$�(S@��x�7����>PA�6N���wv��,�}�J�,�(!nB����@��]5�Pe��×�]���1�N� D%,�t��9���6�6�e}���u���N������(��ɨ/w7��E8|l3҄�˼���HNUc��/��ߏ��!$��k,������5u�Iq���"�2�F�(�D��c-7Kk����9	�����,�N������<'eNH�Rf�ը��?��xq���QEc��%��`�Z℩�}�?�9��Br�l7��=`%�}K��^�7�]���#⧩.������"�m[��O��3ox�s��}
R�@�J�D�C��	��*���#�Ԋ�à8/��`��f��������R��W�^8�o����x�g� ����ի��Rl8M,]W����f>���΢����k��)���@'�� �U,���>d��A��,�Y���
�+;�,����<���%����g�cT���8ͣ�/��d[�c��XR��_��k䪑��T�/�1�/լ6XՐ~3�E7�¢�����ru͓ϡ:[Z�%� ���	�SWp*:��C-�펵��j��ů��S³�MY�0�v���'�Tp0/ kJfw{�c Z��� �v��)���h�To�����*?A���4����5�M�EEw�o"�풵���T��,[2�.e�nJ9F��p���&��-��)�jPI����|�)��|�e-��'������hx�ّ�!"ɽ�O��G�C�mOuGѽ�$�i��*��)�Z���v���9)��}�Ȁ�1D�/{�4�17IU�2ń呰{}ǥ�#���)!5�k�� ��c_��yF`�[��?�����SQĪ�����r�)�}$C@Mxn�:�^i��U8<�������oE��ڪ��B8 ����/0��7PR]��h�j�Z
&j��|HN1f��������ס�k~�JIۨ�
�
��¾HA�L_p�rG�����S6<1���X�_�O���cI/��Z�r����V��G,V�Z���m�r�vFvl2�'�<ܜ<��o��P�%T��#a�lrv�M@o��R9%���O@?�����Y��}G|�Ai|I�����I��d��+v��Ɉ�a���V̰�/�����;z���A�{Ӡ��w�4����1��-$��A�ʭ�0��l�^�W��~�8+�`���n�4dZ���9ʠ��o����9H��G��J.��@���ז��5�Q��)���n�o�3�.l��I�"�YX��z�D�q}�2��ֶ�&2D���_��D��E6��q�[��z��N�fR�.�n��nܑ��,h@�A��Հ�t3o�ɲ�����;�.��Z�'
�,�=󉽈�I�y�]}�z����(���{kM���m�ֹ��'�у��ͩʫ�{�ȽO��\i���Ç)�r��v�V(��A�颿�m���������f�v��Oߴ?��t�]�,�_�ֈ�o2�;�Q�c�������6�z'Y ���[�*�r��olB��{�t��B���8��N�ί��+�9��<ۣu^2�#]���{G[��!�: 4%B}靍�G��z^��d�>p�����@�3�\p�7s�v���xz������ͦCzC�����=�XZϴ/"|[�dF�v,�t���عF_�_��L��n�if��5�2ު��C6����s�ħgQm�nm��)$�e�t��g��A���у���^�$Q�"��;C�ۍ�{M-�w��_�=��4�,ul {�8r��5�?
���{Ԓ��͍�;?C8"�>Ÿ����R��꿯K,}�<4!SDV�`�#�:4vIc%�O�
Q,s;&d雭��SL�Xi�ö���8vF�6g�=���I@��l+���/���T����4�'��.�� \�	If	�|6ç�Ȏ�F����XG�`���/�Z15�0{�:��UX�[�e?r�JewZ���@���3�_��2<�n�S{��m6�Af�	E����ߥ�^�C;c|tRT/鴟�q>���P�q��t�Z��z�XL��c�غe�vɣ�RZc�f᜛�)d2�p�Q׏� W�B���5K|��#�L���F*������|kKj��N!���n�&=�`��X��oF��v,,�����mN�/�Q��dH&����B����=|T�.)�9Bf���S�0U]	(H!�v73�E�߭9�G�_k�Z���X�0lU��
�L��}�K����6_���E���6�~D�c�ye�tf���p�P���+n��Wj
߶�к'ac��qλPC��� �?��,�S�X ��Ai'��C>Vu�8�K��z/�%��8𵫅�nw�EW�3��f�9�IP�$���Go�/�m{o�����F}�g0�)�k�c�åLEP��GW4�;ry�D+S�
��7e��8_��b�Ry����4{�_k_��{�B
����z���J�l0�]���-|/��x~?A�;�^��~�(	�F�z���G62�rͦ��;��g̭���VN��/��h�o&�d�^��.rz�eo���g٤sM�C�2ή+Y��[J���t(��=�)y���*w�PݮIMQ������j�������
Z����$�dLL|�[��*0�I��C�/��Yܚx_R��kv���}��h�A['�F������0���h������Z+���������4�޹�P��t�:d�:d)׭�r�c����{r��X�E`���85�gdI�����W�p�p|��ʹx����@*���,R��;jb��ZdL��Y��޴C��a�;�B��
�I�	�TO���>��ߩ���bY���mZ=��	~�PdˇX���4s�ڼ�w��{��X��f1���һ9o�3��K�岨U�
��T�� w��Qv�dg�.'59w������������:n��y�jA|<�fg�)o��W�ʙ�.7�*�j�.j*&|d�w���Yb�R��tF�s�o��Ů[3"��Cv�_}����3�X	a}�C�]��� Ï�+��(�|�����{#i��]����g�.7��i��^i�	�@Jiwf��O����n&n��L�]��hn�
�z�`��#>����k�ciI�	:��-��9�(|3}'�����W`�~m��_����� �� DS�5ڣ�;�ö�(뽅��׋��}�vYHv`��n�
Pu�[�Yr
�g%FF�T�{O�����@�+�������R7ǁ(���_�C3p��>T��t�P۞�إ��Gc.�I����l,��a�z�"��A�R�Oضv�|{��B&J`���O��K��KN�������8�� �t�q���\���U��K�Y�AF�?�js[=��-}���Ne.T�?�q�i7��xEZv*͒7	�'A29�c�:m�#�#�)�vlշ����ii�&c���"��M2��@� i�,�3�T˯���*3^�wJ�ė�[XT����'G�M��C_��wk����%u�{_�mP�r-i�!`l�k�|�s� �HK�  H�o����������u��w-�ӬE�3ya׆�z��^&��,��U���6�©�"�m�/�Z���L�nSE&���~�ʏ�g/0���)�-0�s����Uʶ�އ��aTf�ȋ�9 ��J�A�ݸ�%d�Rt��S�"n.M�a_�R��B�i��(�GG�~����n.�Y���YmZB0�@�����О7�a2�Oȕ�ّ̅��Q$�+���%�8�6a��|\�X��^��K�hՌ�s����8dI�F�>�DmW�d����^7o�41.1nf�v�TJZ���>��Mf�H�I�Y�@�|2N7Zp�I� 
_�>�2�a�d}�!_/�B��:]�<��վ�W2B��.I�{�
���9X~��j��AWF}c���uw��p��1�Db���9���eb9}a�6���l�<�j'!'#W� �l�U'��A?Ԇ�>L���P�|k�~��b/&���I���g�lZ�-��yw�:���`�T������{a���K��g�'���o�uMCa��\��i��C 
����x�J����a��wȍ��i���.�;��	בi?��
������_qњF��m���^�\Np��ثu����D߷}�-22�K��	�*���'����ђ�4XVw/Ŝ"r�[����Y�tu+�W��|��o%���ӱS���j��(��X�Eu��1!���m�W��Af�f7��,���&�[oz�W��L�o��g���+ߠH�R��/����䅰o_�s�����0�q�V1-����s竿��z�p �[�3D퐥G!���k�P�v��n>k�����1Q�.��QCԖ�a�Z�#��~U�R)���Iz�F'=�/{C-)����}'���:�m�؂d�f���&
A�l�G�u��i�M��U"8^�y��N����Md%C�g �G�
��E�V����*�Dt�H(��ɞP	�l�Z��K�4��x	]92����))H�3�W��*g竽�=�dO�������V�,�م��3z�;��$8"y��_v�v��%��cv �gsr`���/�sk�"����E�����i��Wv�A��Ӟ<_�#��_D�mӵ�oǣZs$9�9�qcW��OZy���~wiae���D�4��MLҍ��Ѧf����3b�&�oj�^j��kt}U�ؖ�3�ݦ�Q˷�)��P�NN�g\�����oTE3��%��d3M������tᙓq���|�����gY��%�Q���N�����q���j,�H���us���,�	�4����k���3
T�p�����/@�)�i�V��4L����0�ȱ���4��ɹ�7Ebvsz��J^R���/���IHp&Sy��"�f�Uj,�T$_��1�P���X*����#dBl�	�]ʬ�אez�3���_��(I!��YT9�
� 	�V������ ,0籖I�q�\0QF�E���H�q(e�u���9�8��_I�N����H����SE6m#����?{߳W7{e*��V��tk��R6���<�ow!<�,�8��L���[6�Z⇆�OH� c�n�L��[�CZ�w�Y�Z�2�%T9?�h�෬�3�od�������Q��T�^�p��:���������t0 `�j�fCtA�x��Ĳ27�f�%ɠ�n$�c�����;��0� �@qo�#~]��0��
�G9r���:���	�;��~�b
'Y{r)	=ӫ1Ş�]����k���X���^kw��� kn���$�$������k&�2K��.��	�@�U�=2h&
��Tϕ�nf�u��Rc%;�^[��Hz����F�����VWKi�%�y@�DrH�?��LP�4u2k�^��������a�r�\�����~�K�dF��)�%���e�떯f���tZOi��U�>�
�Ua��\暈�Q��@�ݧ��L�ZE���yaSн[CS��]2���a�O�B�e`7=���=Ɣ}ՙ��".� �v�U�KF�ս�W���&R��,���%_�U��6:���'e\��*l��]�7�����@m��7{S�k��c�y�o.�N��/4a��&@�4뷃�9��Ӻ�V؏V��K�{���5qY|Ҕ8{�Z]+3Lr�7L�"3���������-Kꗖ �/sa":ÈA�՞�(�8�xگ�oD�$���z#v{{Sba��:P�a�@p��#�v̆�E�l��y��6h�-�oQ�08*N?���d픉�b�"!����3\Mɫ1R����x��D��8�q���w����o����k�/�Ю�55��֧RϾ��`�������Iʖ�lHgf��}�5ϝcs
��ۣd#�
%A��hisgj��󫘔�ڳ��ƒK���ʓ��@f�nm43��\X��γ�w�Q@�j^|�+�u��5$&;�!�1/�b[���y�]bE��~���w�O5
�D9B�i�����f 1����/KJZ���w.,�(�	?��J�����Jb!yv'���;Å�(���Ψqѻ&�>�W��ʍ��YEEl�2��i��;O��S$���gR����b/�~6�S>�}&|o�%���� �_%a\I6�N��&I����O�U��A%�w��f�W�, �wˀk�g�jy:����ԯ�	�A�`�,���Q����>%lhp�5�����~�<1�����G�B�+��r8f�.]��!�B�q���!�,���E�j?m�h���q��!T7�?jd�ճe@��;9Pe����pw/���/�b]��TLO߿Q������K�&���X�rfJ���)a�읍?/����"��,+��T��J��)��+�WH �C(���n��gpN�C��+2R+�(��M<|;��@:ئ�������y�m �zF�%�Ff ��Ϲl��h:��ì��@���_�mޏ����)��߼&�z�O����rHt�k��u3�N��V�-6�� e���ʤY]�cxJm1l]b��j���;4��UNiB��;�n���c��"�WM���f���͇Z�_��w�B5�'Y~лZ���I֓��'�O�@K���:+�&ltr}�r���%�H��Q������,���g�ł����t-$P��IP��mڐ�0���<XTΎ�>l�q��8��g^���\\<k	Z7�����R>6��hWN⊶?�p�9i�䷚Ge)�K~����4I�z��7�ow��5�k�H��Q�2U�	���-�v����"��%�����Р�tK���l�Q2≮~�F:�-4�
�$`�V�*�?ܸ��%W,���D����
�i3���i���{z�vıO,`���s��.G
��`�6�����⥫X_y�����Ԑ���d�*���}AOV�t�����4l�?J�h,�Y�č��1yk�'��q"I�ii�(�`"Q���$�R��覆��:��t�vO-��ysi2:�������+����@�fӛ^�������!�mH����/���?��x�,��ͣYg�\JV��B�D�ۃ�8d0Ŏ��@4��(K3ס�ixC�u ����o�E�l��e�h������	��)��ވ|xP��='J%�3�����k�!��K=�W�_6S�`��\��� �՗�?h4t�yk�s�.6���7�r��ހ��;ǎgN�K  @��$�z.��d%=��ҏjҸ�&�&o%y����]@0S@���)Uj�voE?d�y�;Iy;�pH[u�?��� � i����:�t�z� cW�y������Z�3���S���/���t.����.�J��t�G��*�j���Y����/�G�>-�%���1]w��]Vi	����7�p��ap�ŗ��:��x�w��ԓ9�����E��v�R��,���d:ҁ�$���O��K���5)�����?���.���Լ���@c��';.�E�;��r������P`�q"��L6��z��&��k�L�g,�ɮ��]X��u���U���b��7�݉7p�P�1�;����5��WBؾ�(���w;��}�z��Z�u=���M�eHw]�݄��[��З�κ��!k�C���y`=�P��	[�x��16mIq]���ž]D@ u_D�_j,���i�m�X�(�b�]�>���5��j��e�;t���(mj7Gy`�@�ӝ�j�۹Y{����'�����)�����''��R� �3Z*(�0���q��>
����>��9�i��!���Է�}�*���"� �I־�=��Iߏ��;��P��;��Э�.�W�!��ީx��ɮ>}�4�3X�i�~%G�a:blU��:L���|]d��9�:���d�aI�<u�\�-�����X��V*���/�o_V�a����O�Z���y���[
*��B��P>T&��߄�K�#8�f�Ї�+b���������x�����8 s�4{�c���ӱ�L�,���Z�v-�6���
i.2d���!�_��i���oG�g���>a�'�
5���� ��s0KY��K�j�����DJ�*`�^(h�4<�L�;)��h-�;���^�Iß�u�>���|�>�J,�rc�~X؍���k��x�s���m���VA�7�0��kHz�ka�<�sNm�R���C)���r���HMK�V=�
1�;��܏���#���/\_1�>&DQ��a
��]��UK�1���%�e'T�/�����k�P�Vye���MXc:?�I2���{��N�f��A?�/��'�a܉��*��&�ۋ��᥇ӌ����)&Yk�`47�G�I��X�/���dT����˵���XC��O] �ҁ������n^V3�'��)/xX�=�~ �R��ppA^ + CP+o$��C�]_u�\��^��|���%���v�~��M-6h�ɞ�詒\�ŵE)Ƭ�p�F[��F�mR;�y���K��[��E\4���F�KN�����f���ا�]~�3�Pކ_�>�PvsP�Q�I�7�H�����%���'��w�~0,�,�Q�m}�T��+J���r��B��!K�C�?߫ 3 ���bi3�gL�K�~S���c�| a޻��g`C�U��q?(�m��F�<nX�&���V%�R:��Q����� ��ݥl�S[;�k �2$�n���E�L���[�I-\|P�7�h�( S�~��~,��냄1��8~Ӌ����( �4U�R��0��EM t�|h�@������*���g��Q�1l]�e�Գz�N@FK�J83b�܍��h��x<�i�v��kW�lv�t�ܨ
m�m���{��,��E7�s��]�v�x�����]���2F���m.��#��Ғ˹����ߡ��T����U�h���V��Z=��O��yڅFiW�C�56W�>�ÿA'AI_���x�B:D���.�����l�o�dk��ꗚ�%�Ʀ
#�$H��mQ?$�	�������1�0.�R����>S���C���5�a����O#%U���i%B�Ͼ��k�ş�W_�	���K=�o�V,{?A���@����d扃��#���k��5��|F��{�=g� �0,���t�e�IB�d��G��v
��l��`�ۜO��sX����D�K3��6�~��h󩭈�����Gj��W��p,�S���1#R���
)z�d1�֠��L�M�R��2�_�\�����aj�\)S�~�o�� ��D����ڴ8$O�	6�'�8����Ɂ9 wtߝC��p@ߚ�545���������E�C4����uw�.�b���!�酪a3���Q���d�\��qt�_�J��@�9���>Bu֩"�ǖ��%DZ?�I���������)Ϛg.���.Ų\��
*�x��xwE��wt�ͅ5�O ��Q5C@��U{��%���ڸ��7��KT}��v��!�`���@6��58���3����j�T�/	;��v��4~��˲]w6������Os� �;�xT�/鏒6��6�g��N�-��9#�NŜ�]c��L��
O)�N��E�Zx�E�B6���A��Ĕ�U�)�{s�p��\1GJh�5�c+�@�
��w?�����v�z����="�� �5H� 	k����&��j�]��Z����T0�O��x8�6��������we���D}�j���f�ZӀ��O|�K.k�nc��X�mU>HOKJ�.����6�tN{�Tv��q=� C5pW���#}.�c5 �p&�k[$�c	1�w��z^$�r��P^�, �ͻׅT��O���]t/ J{�T�*2�÷�V���x�<��ޕB�3�.Di�����u��w�X���F]:�&��Dp����h��Ȧ}1ߪt�M�H�a�Q��/ܶ+�ё��N��-@pt�V���o+�����.z�1pa���CW��,�}��o��p���׍(ƏF��~�ŋT�z@]��Un��.�,z�-.�AF�Rך�;kT��5�d2�"�O [�xn"B�_�$2�zS|����Vp��,�$�k�g��/�a>i	:�ua��5E��"�ๆ4� �J��^�:���u��;g'}�+�V`�G�����|�ׇ��[�n���]��x�!%Y~�J$ӆ��v{��`�h�lyRU�(��߮�%{�úf�X?�0ٚ�7 vѣj��'��YT��B݇{�?5������+PP�*����*�Gj�_0�MPO�n�K+�ܿ?� �u9�GN8a�d���N�����S��S�������L��D{�ޅ�x2�=+�ae��B��|��:�u�=h�)/�ڟ"ώ��V����Q�$�]
��F�G�cՒ��`�"B��|��Շ�Kܜ�}%̞�G}?�T����,^�f�yʺ�KXȍ��7bW�߾iװ����Q��`��|��Nw4H��6��m�.������H��ou[PkxC]d�Y�5@`�Is���PF��A8�yO����x#����e1���q����w_srU��W($�<�JՊ�
�+�y�T��ajS~2{oV���TZ�d�_&���|EU�����T�f����U@����z���V�/�n$9�)S�J���f�c��kz�5�#]�Gȉ/;���9p����h�&�1��v�ik6��C��T����.B��E�,�;s!�1�-��6R��n�]
��w�[�N���5�ӕ�%�g�X���8?�ufv	�����_@L僡�6?j=�� w���Ir���\r��9����GJ�����m�~ׯa&���c�W19g7�}w�Vc~L�~��nA2Exܧ�7�-�5nR&A6r��2[w��w�}�S��z�yՆy\tȟ���SxG�H���=��/b����91����Q�f5��<Ey��Ne%%'&�Hݎa%>�J+�raQ~� I��JʪB���(�����x�[ŕiTUU��lc��>$����;6[�����d�2�'�'�y+�=��jzjjUm����ЯG�R:�'ܾ(��gzg��3B1�f�h)q���7��˥��Cђ2-J<�Xn��e�Sb��'V-����in{���*���j��%!Zn.������5�O��0�;�U���x�T�4`@~i'�\�E�����iJ�<�z�ڎg/[L��.<��t3�U#_��ѿ���&��;zx���e�u}~T�p�9��Hʨ�����a�C�d��%��_�'�+<
�8
���cMRj�]G��m�y)mٴ�_�ߪͨ��;���K�>��b�UȤNl�i�<`�k������X���l�Y��ҹ��`3;['�`{;���uP�L��?�9=��Q`��jH�+F��D�^M�v�yq)T'ey��[�L���u����3x�(.%���՘�����V�y/��_�^�����;m�*�{*��p�ø�yǣ ����n�4j��)O2Ne� l��9^����>'�w3V�5G?E�Vm�5l����Uv�,z�
y�r�M{O�i�h��{�����9����1{��R��6a�Ռ*���'�o�4i�$��^�v�V_'}&[�P�[�ã?+���$Ûؘ�L';�]���&I\S�%m�����b��y�	=u��Y;@;f%�!��;M�B�Vs�v����V��xV��O��;]���׿.�����g��;t�p +�'8�C�k�(o�!�)З;�z���[-�X�6Ɖ��i�rsaQ�-Q�����aˣ��_�ݸ+��˦U'+Ob��N���)t���<�ƙ x���,�4+l�]}k!\�Q}�Dq0�궧�K�P�Z�΍�1��xc�iS��v��+����xX9 -}.�j����?�� � �o�{]Z��5~��$��x`@��W��N�?��2W�%��GSF���NT0eN��w���TxݭXQܗ�S���Q�@�4V3�2�+��+�j)����W�t��h���4��8��AfE�Sވ}&X��Tbc
{{�$̽?��C�:����x����@G����2Sށ�U�Xi)}�$�����CQ7�K��-f�M[�UC��A׊J�C�S�S�m�0H���������ߟ��E�����%;Į� ��®��yuǪsjq%53a�#���&���. >�[����;�k&~�<~��8�����<��nY��n&�׉�'���N��q#�R�.杋������B�ki MY� N�V ��0fJ����6��[W{�S}}�W�X?��Y�k��z*#�< %9N��
ѯJ�CUa}�@v1s?�P�hU���� >*���ě���&^�U��~�3��r֥�ԙ��� �B/1�?j>����_.eK.���V� ���>�O�"���Ñ�U�R#��Xnϴ+zU6N�)�m��ɖ���� �N�~�;�Bd�{y٪*�+mL�է�|uB¤(�-��Y~�֞�&���g� ��Z��y���;�\�|M�����&����ԥ,�4}���q .�[�RK�:@��y@2��Z	���,]�Z������_~dj݅d�8��jߡ|��4���o�xA���C��U�-Ȯy6\@Q��R���|��aӖ��B�kݲ@3^����J��x�~d_�>�k\-^�U�^�J��o�|9U��$��w���ɔ�����[
w���}� �T;�GfM$���07M���~�E�k�B�'�]��\^��3�ϰ�uOƏ7�V/7uqܙ�ö;�[%�, ���ʟ���(�u�%m�;N�L|x!V�5��)������ֲ���u���M
�yI$�0�_u=Vm���_seک������r��`ՆU������m��i�n���tcy]��{7��l�����7���|r��QNN�؄�4\�xCM��g?V�}��1��a�O�m�;�n�iz^�u4�q�Tyh��e�t�"�=���0 �#�ڀ��N�P��+a��vG�\�~�%L�u�&�[�EF2��o��~;��)���.2����+���<�q�}�I�i�bK�L��5к7Q��%<�z��A*����4��4U��|��a��9k�NӬ�.��H�X"ŉE�(�����PZΡ� �'!�ko1/5j1�ک��YP��<��D4vyc�H��1]���bk���]cO7���;�zpПg9�M��Wo԰E8��H�e�'$D��W�����K�z)���G���j�iI��G��^b���������1w���@��;�y.C�O0�v�;���h�n�Qk�a`fs�꯭��Db/�W�"�M�?������议=�	�1�z��a�s�g�L�'7Г��G#��s��aI@��`'���/��]�]���vfƝ���1x ��P���<͵�3�B\]��u����6���s�	�rb��ۤ�������U��'#����X���s�)���>��y������ۮ��V����h \4Z��E�&	��[�Z��K����#��c̟ޞ�w����J�_O�fF�h��j�c���7w��"��]x<��jҜ��'Y5M0 �sMO%	������e����kT�AUx��o����}�$�b���N�`��co��xD���?�	��_�|j������7ޣԐ�M����b�@�?��%r�j�M����hbZ'{�\��d���O����F�OG�y���8y)�O�5?�g��z�0L3����iݹ���˝`C婙��j��_�ɫ��ټ����{��n�`=���:�����{�ࡖ�jJ��ˁͿ�v��캆�h�6��]AlU��V�Sߖv_������� �p`T���M���|-�w1кa�dd3�f����/q��7��Pe��)8
�I��OG=�Y0RQ��P���Х$��U�4sF"�.��=z��;�̈́����ۅ�30�c��?ܽݜ�5y�ձ��C���#U���	�����qm�ډb�Q{�Ȝ���w�v����RAyb#�>�6Mh���6C8|t8p-�0�d/G̞�Ɵ\�$X���h���>�~[���
�]��&،y���GU�xFT@Q
�d���p�A6	��)���_�a3ح@�;��1�>*�j��M�Q\�t$�G	ss���n��Qu{��#��?c��^3�;�Ȳ4Ҝ�,ڣMʕ�V�ݩ�����פ����nnD��o|��)<{Q%��{��e�i�i1V��c�����䕮�U��z3��]��S�ƢA��J��S��@���m�s�B�Q�f1&����J�1���Lv�֓=}ڥ5L��3�u��Wi�hR��;ZԬ_���0b]M|�����n�_�����j���D�H?�^�Q�N�m`�^^%%�����?��9/�@�5��n��5��f��Пaj���g��,��w����ש x�[����klщ4�5WdQ�E���;��( ����l1m�=��/���wf��(���x�@�o�� 1�o��NQ����G_�˭��&�8�YVp1(x�KO��.��]���	�m�S����ӿs���y~L1"�<~�~Kc�#��b��W�DH��z��$�#���ּ�cn�V��:���!�g� �:8v����Ӕ?�I-�$+ v��s%߸Π��h�KPL�#l��{�gos�[ױ��!�U�ӈ�G���)]����N �Cu �I��������nB~q���%`'������e�bq�,�&��桮��j�'A^i`���h�ub�%�.�'?!�Pg��#�I��/yacżJ'/nq��/s�
�I<�B�ȝ��[y�?/"�o�;�s%�23�O6�粒�'oH��q" ��EA�������<�����;�`j�_};p��|��a_L��)|�� ;�u���taM�mU�I$�s[��D,�03aKt���f
*B�kE���?����+���b^�/����*4I�HHšH���pSE���#�����ͅ��m�����j ~�ݎv�rEt�#���x�W�p���ߓ�!d����3-�0ET�Sj���_]�4�|`(teL�hu���4q+���K��̎����3��_���w>e|	lX1r�=];v�A���zo����b[O��?s���K#�ڞ,���`,o��}Q�H%S4Bq\�eS��	Y:�jGL$��D�c�"�x'H�ua�4�_Uk��cmg �.�a�Ɋ6��8��T
B��}�]�	�Q��	T��\�PͲ�'�"�B�f�KX	<:&��㦍9�a�9�]M����m��y��+���Ҵ0��<Y��T�M�0�K���Y��Aj�4kg��;M��7�+Y-�Y5x�>'��5�����B��P_�������b�^ƽsVM��TSn<N:@@�<�U���,̲Z,��n�{t�k��P>`�9Pq�|>'/r�W$Ϲ�F5 PԸ�C��8�Я��nF-�CrW1]UYM�q�jG���gGT�"iD�w-B� K-���gW׆�D�hE8B�̗��N�9K6�jWۀ씚�����\q��RWخ�jyD�2��O?����m�n��E�@U)<�:|w���JH�HϢ�@�X(@Pf�v4�vy�u��j�����:���W�W��+v|�3jE��>�5fPh�M�1�?_��o���9
>�;�+N���?�;��ݣ�'&����������V�4�ʓǿ�ϭ�0�m�s��>	�}/ H���G�c����[�:i��ve'/бOax�f&8��Hd�L�u�-9�qP���e���Y��2T�!9=�z����R�x�(>D_��H	̫~Q(�W�4�?k�V��Q;$0���#����v~$�X�~�u"u� �6�O�PRӥ!�2`��Zpx��T[�� ���+����a@��K��c��DL*^�]]�Z�m��!M�g9�2<S��LO3��j������_�b�hO˟Յ�J�����ޖ9��@^�T�@&��uD+���O������ �ۑcX���@����`�,�)����b�@�ؓ5hgM ���xX\���7#ʓ�K��3g@��q��)j����|�RJ�!c6�c	ةuL�ο�J1�{��؋A�Ӽ�ߋ�eIuR	�I����gT"H3#�=�!;���� G��*����_�_�/�d�����?o�5��j��J~�9�j�./��2�9���&bA�X��z"���.�{h�ۅR]r9{�_i"���}�J�۰#�����#Ӈ��	��Z�����)����+.!Ƴ8h'hw��VE �)DD��~�Q������&d���@}c44���y�!B2���Xr���Tp��z����!K�DKef�w����:.��k���*"!R
J����H�R��0���(5�*�"�1����H3��59������������Z׺ֵ��g�1��j�`g�4��$��*d_�v�+�M���S�_���&���,)���\��������5�C�Jw���v��כ�yT�U�`��{�&h�a9oP��v8<��_Y�O���@+�wӤ������숕0o��iX�he��f��M�?^�$x�"��	S�An������?��3/ѐ���G�0HȨ�
=�'�̛. ۬N#�n�j�¹�AH��q\���!th'_ǃ�K�OE�g�Q* �j���:��t�^`��]a�+�m���MD�A��l�q4V���}����������j���+��7�����46D�hA٦���U����*W耤���.���[{^�BG�Ô�$�>�1WU�Y<C�h#꣤�S��uf�4��Ƀ��6p�����2����hd�yf} �6�hy�YHR�ۏ��s4�
mH�n֤RP���6�[��,/���D�y�S�{�2�}�����2�Ě�e��D&�ȅ6rīn�yKb]N�D�D\֚�60G�cYn	&k��)�	p�ι���l��ڿZY�,�`�`jBa��חn��WR߁����&T��H�!6���@��4��]s��\��S�)4{!hS���v˾�"�����GBS�A��-��W��?%��1B�02�`Y��{v�/�5SQo~�����_Ǌ;�5�@2�G������W���ͬ�='��P	M�_uo`�W��u��4�S~�*Z'L�OMR��_:�\��3]Gl���r��O��ǌp�l�E�k�A��*���>�*��Y���\F}�t=PgC�~V�++0ph}B�o�ľ��y��?��*����3�G9���[*a�\t.ߦk��0w��@QE�}��3������a}��h%��o-#v� �e(�%���D~���M�n9�A���DO?Jt�tV��wl����O���f>���j�u�Q[�`o��	�J\[��C�?�y�ݠ�w���"�L_xS;Y��B^<h�g�s�E�)t%����Т�Y���d����W^��+��=�$� g�uɮz�鵻�go��y�Ys�&|V�\B'sx��܏MR����j�䩩'�g��K?kTR��g�7ʆ����1�?���݀�Z]�ow fzM�jwt�XfaYz/!3��̪7�z�H4��/	D��g�ӛ�#5^yʭ������}2���������,���Z'�$ѡ����Jy8S���6V�7Kr���_�_q��a8�o[T���Y�vz��ThA��o�8�B��wQV}��R���M9�s�<+6�d���ݗ����8)��[�fc���|���~s_
?�q�Nw~�T˘�&R5�F{707���m���֕lPzk�[r�N���F�C�`���6�Cޥ�S�-1O��2��B;���*ɩ�8�@x�6����@h�I��F}YL�	���{�����M֞q���ER�&/�]���Guƻ�c��U��9V"R�x�ӡ9e���-RX��=�4�lmU��G��K��T�35�8^7�q[����dO���M|�J����P/*�9Ս���v��"��y�&�f_��f<;ɉ��>��c�|j��b�<ٳ�Z��@ؾ�aW` j�t�|w��
��B��+�#��L����jsq�\ZL;_��hf�^���'�����Sh�ȱ�!lB4�������%�_�w_k[0P�A��7�L��3/;h͙M�4�p�����+�^_�����j:����]�o�Xo��e��d���z���Y��x�
��AYl��=���4�VE��7�0�-��^��Y�GUH�9Y�&��ճۨ��p"q'���M&=L�>31��!y`p��0b"�aH@W��,me}��[y��HZ:�=�C�j�;�����n��<Ͽo��:Iئ;I\Y}V-��>-Y�F�'o�{�Z@�P��1ʝ��Z�{�ٔ��>R<�]4=���@�`q�$� ������][�.��r��|��Ķ�����UDAQ�͑d�9�<M22��9�x�|�.��������~Bs���;�+4���P���
�Ƽo�i�!���{]i��V��Q��
l26�_��$�kw�9v%���ڇ�C�����TTt�ӻ)4�$��S���oWΩ�� 7��qgv�ͩӔ�)�@+S�[+ۭ��k2|�0�kӷ0M���)%�s�gM<~��n���32��/��nQ�_<z�!�5]��o�G�ƴ���%:�n�������3���=��w���#��l_4R��X�	'9�&�3,��4X�.q��cN�����R����X��О����\��h2tgܠ�i׫̈́��v��)3��8�"�z͸�{�y��'�<i	ƭU
�V�*Vj9yq��}I���	���lL��n\�S�k��0^�
���i��xP���%���@We�h�����j����Q|�x>$�N���Z�w')�
L���G����\�
�Oٙ�!|�3��`�u�X\{�h������m�� ER��kz?���~�R[��2��N|f�頄x�`�����B�ϜAn4\ʠH�t�`RЂz�"M
q����N�s?�S���}����<�dq��`��(?{����?��{+ʻ�����ؔ��ZB�7���]͞�j��~!�����w���h���w��dK�Y� *4�z�U�جT�%�Z���_���
�A����`��s�o��q����,w��W��4�9f%�Ŷ��DPx+ͨ�:�r!��#�v3������,��Y⢈Ec-TH��^���	��I<��'�gz�t��h��p���͍����;�׭��&Wʦ�3,��j��w�JTr�<���˞�!���iMm���R�����ߖ]�ﶍ~z�E����nx9�����)�S�Cr��>��ǜ�Z9���s�ZfS	N���S�P��a�zjm|*�װ^dv���9��x�9�9��/x�U�	"�ľ�&��K���&��y�T�	Gڮ��b���~��u��Y*)�ܨ�w�����K���S%ߎ^2�gsG�� ���v�Sle;ت6��M~VhY��Pr!F�ˮA�/�3h�W��hiT��I��o��$�]:�CH�v�����91~Y�K���#ô�X�_dCz�-����#�M���R�r�ގ�W{�j�9�&5����;���jR7$�#�ʞ�.|�I�j^�������ņȔ�l��mE�Mo��G}������Y�쾠��1~�
�F��O4�JyJ��[1�CĠ%�fq1�u�R-E6?{L���6TaQ¤��^�T����@B�;p�o�5��ߍ&|��{qw=�a�W��;ǔ��26J�!U�Cb�Wk҃�W�j�� G��?:�3}�Y��nJ6�yQ�BU�?F��J��Ƣ�w`�OQ��Sz)�2vfojj����}	 	fi�b�C�9�e�]t����՝��PNְ���{<��h��?���|��|}���{(���� fJz��M{k��h�[�p��i��H�r�X�Mܒ�_ ��)4>��P�S�)k+f�0Z^�)Xܼ!1�\)���|���6}Wԣ%���BQ��G^m���� ��Ge	�t�wb���/{��SԤ�%w+�/7Ɇ603Ngi�z	������//�m�����uW��.�=ϐa�����t�����b�Cb^�;��K�.�Y�ֺ��ɬ?M��"%���~7��a���c�G�s�^�G�ݝ�n������i�a������6O�]R@���Ϣ��U�i?��������[h��e{��x�c�0�+�S?���'� /���06*mą͜ـ[�! ��n��'BxFV�����fxQ�W��{
��Nxf:�����g �;�\�����[��.FӪ�RW���v�'}ʕ
�
w��;j��#%��y2Vm��	��)��lN��?g���r�u�e\����R#����ڇ�c��2��N�>r`bb��G�����0%\�]Q.��u��G[��O��v��/���k��N�ܺI<�]%�	�_���jV�霪 ~>'e��fdX{C�K�ӺjD����yx�ޤV���
���,��ܺo�����t�y���V�d�����Jy	�	!p��Z��/��^6����R�V�����2���u��qq�"���?�}[�ﯲ{�.�ȱ3i�P�g7�ؤ�� ��c�h�:Y����ˏ|�kht�;�h�UeL�#4�V�vwOd"S%/�U|{@�<^�՟]O\���M�҆=�s�Y�_��30O�J�ϩT.�վe��i�dn�
��T6���j��K��M>��yK�Ն��l|Qf�Z�j?Ea�)�=е���kR�@wS4A�v֙��0����� ��?���2�����C�m�&t��o9���N�A"	�ϼ�^��l;	ʽ�M�k�c�rU��|���$��&|̵�c@ՅI�\h�;#=��N�qU6��~�e���|;B���|�Eo-a��w=�
��
I�"�T=�X|�����D//�~í���}I����R�Q�M�g��w�mA�/�����-��4������؞�ӽ�:͞CR~��e�[ʠ*͑a��EH
r&�t����3��ө����0���o��
>��ŕA'��T�jO���>�η�]���U��m<�_ZEB���n�Kܴ�"�� �aﴫ&�jJ��މ�v�l���ݙ��x�Y�+�6s!��>7�k���^��}E������+������[-�t4��tQ~G�GuQ5b@���Y�����;UƮ�ɹJ�y�����Ի�Ei�Ѹ��v�#�3��z�ȧ���0$k\CIܒ���1*�W�hדF�g�hrq�N	� /��:��`5�=�CT���!��Q�I��X�O�LSY�����Zhtr�'(���I��9�g�T�:|.�(}.�tJ��N��祖�g*⩟,~��gMn���i*��a��~8j�u��t膁���%�;�ZQ���>���s�>��TY�ʼ�v-6M�M�5��t{;��=�ؽ���>��aH��$GiZ�TV�C���KC^��y�2H��ܯW�"H�3�gQ[�!��/9��TL�|X1��H�=���9}�8\�ޒ�,Rya�����b4n.�	�CŃs�;����>s�-�@�^���2��v��YN�.�{d�|��m
+l7m��{�ᘍ&�j���Ǌ�;)q1<���;wA,*Q�%������bȻ'I/��^���w�L�@� 9�6Q%�͔����Џ�Nw߿3��\���]������}�w��K�!�>Γf:o`N���'D15I���,t���-)`6i��B'���ǳ>���?w�ն+lW򄮫�&�1���Q�	�3�p���;9S�m��M����mր�'SAE�<*:���$%� ���8����m_[��(˟�>û;q�	{�d��%&�����O0�#�Dpۋd%e�YR��S�Qd�}�8ja�qLm�|���L��Q3L2k+�\Ko����R�=�U�c�A�e����lġow~TT�E�㾘Fx]3�_nVd��PHx���V����'U���$�4E���0����]Q�A!�5}\L^�n�@��������a}�ϨN�p�}����	]� +J�\}����m*�����d�L:�:�)/Q�12��|�s�'���g�s�7��E��c�=���Ϛ��W�}�?-9%���:��T#;��h�zz�_�:K���h"���^�}�7\�5Fn{�x_���J�(e:+�-R�I��e>�a�)5\QU�M��v\��>�[*Ԫ�^ d��T�W�^H�(@~��|+���oe����}�ͱ��xa�؞����c��X4H�*6��T�<�� =Kw�^����|jE1�����gO�@!���_jK�kLD!�jw�Yc�MloM�W��m����s��^x��;�P#�μ^����N��aO��r~���w�K_�8
djB��Sk-�<�=,��~�K��&�vfc��5��U�:�
w�61�5��y'������`������QUO�C�al�/�m&t�G���x�J�+|���`I&eo�Ͻc��H<��ʷ:�H?L�j�NVx%I�|	�jJ�ZK������f�̢t���r��4��64P0ˑ�9l^xq�Lo��\c�HNPn<k�����{����Ť�f"��],q_b:�M��)�
|����a��aVW���qe�]��<�-�S����%���������j�g�
?p��S�ފ��B�+e�7J�?���<_JF�u�c�6Ka��=��$��S��~�.n@Wp%��gNN���*3r��|�Zȵ�1��=���nvK��K�AYbd�A18x��K]��Ix��if�B�p,���w3K� �h��<��3�Rd��A~��Kt�3C�B%x(��X���`�^M|}<+ ���J�(�Zlw��)ͩ�M#��}���y_�P0�9?4�=g��"Ӝ�t�����Q�f�N�l�����ė+K`o4��EW�{�����H�� W��Gd	k��?�CO!���1��zt��ϼ�$�D�����ѡ8����n���Y#S%I��+�+��ysI�JҖ���U�3�;r�
���B{�}X��2%����b䝣Y0�,�M�aLP*�C)��-[$q���[揎��9�]X8G�Ն�w��,��e�k+��ڢ&$Pռ6ۧ{�~C6�>,8�^�_Ϟ���b� �W�)���j��~,t��q���B|��S�V��ҫ��FY}\9A)���'��g���^k�v2My)����`�&�����2A��7�9�*k0)">�&��KY�>�v�n3�'v�<$<����dw1{3�\��_�KQ	4�ޘ��M�ޘ+p�oJB��UJ���8��ɕ����t�JW�GC��p����<��]?E�q�c�'@�Rt�"���H�۱i�D(�N����/U��\[��y�B���֜��Ѳ��8jpb����K���>+��J�箻xlg�^�Ӈ�Q��5��R���EJ	��"�j����o�)Ooq���|LDÈ���˛}ZO��U�f�~(�E���*, 3��6[�o�����/�����a���ͫƦ26�H�}W��6���nD�M\�yt$v c%	�G�I��?Tb+Yb��=�۳Og�[�[���=���C��P�f�u)	0(�a{�G��w"t�?�	�;#�ly���X�~T?�FS0ǁ5c�ώ�Ѵ|����G�(��؛):"e�����+�P�0{�Q�ݯ{)6e	i���'�����s�c�@9�1��UIp�ݮ�+z+�)a���7��e�HӺ��N��VS3A���� ���l�9�H<�n�T(`M�kd��[�mc>J���@�nU)ģ1�D���[�����Qz��?�"�UWq�]Y.���� 6-$̌s�y ��&l�t��'�d��d���*���<�r.\ niT���ރ���{�v/E-_ۜ�|zț�³'��sz�|Zȏ�a�59�ͼ�-ȰV�mY~�������e��d���5�+4���vDTK��6��q���@d��H�wK����w�M��݅jC8h�3o9�/�_��Di��=A���r7�?�~��Q�~����\r�<�T��=*�VbQ�﯇L5���@�y��K������ ��&Q蝥�橡�-�4$�Z���T�}Lp�����;P+Ϗ�<�����{�(Q���t���ק/�k�@��=����v�1s���j!����K�_����,�+1C�g��7���?���{V4�U�����R�rS�����ɅO���Q��$��ӚR�&�ƅK��� �,���q�B�ևbA��%Nv��8"�^����#Wb��r�PL�a�JjII�2��~�y�e�̒�ow���d�0�*�2霯v_��v	�A���+A� ŌNb#,f�W�[���0�ѽ8�;G>�9g�G������,^�I��EZ�i�oYhA�rܑtI��>�7�V8���[��a�D���14�>E��Xd
���Ύ0��Y�ud�yR�6lb~]��t�H7T}��;��f��i�_�2��$1i��/YX�U����8����*��Eٙ, P$�D�˻0����{Svw�Hj3��4��P5}��"3�5��,�U����v�@���)�Em�
��ϒ��VtP����D��8�N�����ށ�~Z�*T�;m��!E�]��ȯE�I�g擟��|��ܴ�'/i@[)��F�S��̳���|�u��S�53��s]V{zgIdU�v�(C�=��*���4^�">��	�P�`�M��[?���},a��T�I*��á���-9�Ê'�\5[��c0�Z\6��!�����C�+��M����܋�`0�v�6�wst�p徥4Yr׌��J�6��m*�[N�B�;l�Ì��P�s��W� 6k�:k�5&&J��mگt�+	�E�S!���{�}�Ͼd�>[^7���������`P��#�PKO�[H~}�@�(!�>ܱ*���f�@~e)l����,�L1�ޛ����y�K!� �0t�ɨP!�fǭ<[k"+p�o�;�է�ln�7�(���xDنތ� ��V�8*�j���9p��Y����q]1 ���aY��qn���%�C�N��(8��f>Λ"��1
��=��Xyw}�G�^�WҔ�fe֓U��Jo�b�^ל�'�cy�>޽�cF[^��]ScP�Ǔ�Z�O�I�"E=�̯�~���.�רf#��k���xT�7���BRdq_N����/#���o����W���(�1m�Z��o^�~��� �Op!5�5��6r��=��$\�J݋���^=IshY�P���(�N����/���5�C@�����
�9����s3-�H-|���4�N��.­�ਪ�w�)H�/ ΃�߼�����ٛ��_��q�q�{�Wr !x�.>:���/��x<`;�TQUB�\���'�}��*��C�������!�S!'��v�cve�}��yb�[l��bK8}k`Ʒκ3�n��j�9z��Hҧ=Q�H0��7��Q�������MӣMT%*�����0w�bV^Y�I��7E��m���iz5N
�绿��[l�Nڋ�F��9�IZf��Ws`�AXkD�	9/�IG ���қ����\1n�}����x��n�1�{�O�
P٫�LF���/'g؅/(C'JRl�>M�B�<d;�(�F�����FO,wj� �>����VR�/�?�E��v�4���@�s�������Un� ˂��� ^��b����6361˿���^V���]��z�JA��t��$��7�5�fSTF��f�޸*h�����5��;�Y�1&��=�/^%��h�*���9׆N�
uޥ�H�WNj�R\�J�-����~��8���r�)n��R�Pi���ߦ)�l�6g�qm!�~_fZ��\Y�)|b�����u���%-湐�d�/� i�$�w (�a"��1�����(�VN��W�ϭ)g�Oz��!_ߟ:t�Y����K��^���#�o�P_�P'�������1m�ؑ ���g��y�����_�X���㘋p�i��ދ��ɔ]�[�Ξ���%P,�A���N�]���lL�;���	�Lb�8�	�	h3"],�g�A2��/V�肞�����#Y9%��Wnϋ���6���ʇ��U8��\10��?�)��	�����S9*�� ����Lȁs�.1�kȊA�ӎ:U�����ٶS�V����P�_(0\Y�qa�i��7H�H�F�"A���۵���@���k�3���	���]���Jl������l�9��̏�p���W]��"S�}[i���oQ&�>z�?vZ�7mmk����'�Bvk_]���.@�aa�ِM��r,���E�f���6*���β�`M�sgQ��n�}Ҝ�{�C4�˙^;���dٽ�M�RN�\;>��F�YH�4��*-G"<��EX����̴ܲ#���M)?���Wa���`V���g�O�(�c�@�,'T��mB}���[?��E�\���;�0
IC�>�����������1�I���?A◿��q,xI���F�@7�<�I�(I�n�|�w�۸�J����id�4}�J��Y���t�m��<'��`��:E̎�'���,����d���-:�����ӎVsa\j[�\���x���jg|GYyc�"�ty��|	�{��8� ��58���'��-4=]�BKVDn4Zm��=���sքɄ����<�%�h�ϐ s[MzX�m������:�XP�V,����4�]�@_����E�o$$=�rP~���qm!���+u>[��)����!5ܛ�ŷ��EVu��f'���˙�S��w���E�@�8��w���m�ڍy��|��st$ �]�f�W��'�����sK�-���k�ީ�I�������J�z��"�4xg�� �`��G<q�l��B�<�9Q~��sVQ��?dXr������w��L�'.T*�MRR�ܿo#���
�`�X��N<QD^+��?|}c݁I��K[Ǐ�7|(�L�B���#�}�T�?��R5}\�b�ô w�x��4�],XX�j�C��r^���{�W�e�q	�3��z�i�J���7��dE}v��"O����7@�����w�0���̯���J^Wi��T�b���*T��!��}st��ީ0fy�q+OLҨa���%Bs�N�~�K_�;�V]vE�u�qɛgP���}C���$���F���&���>��ܲ�@��p���c�y+QZB�����o�z ���)���Fa9d�^�Z��IQ�ñ�/���*��������E��T�`ߩ5����aeD���L�N�m}&B]�/=2���6�u�
��W��}�ʦ����T�/��|�.��+O�{���ή��U��sByA]v�k#�������XW3��+����N��܌̮�:���P!��C��5��a�����v�����N^|���&� ����*�wH�F��p���Cjg�����=�;0�CMs%ghuԑ���bcd����HL����L�œ�LB����v{�����=��G�Wu3{����$��c��1����U��_��<	��6�^��a�G���5����W�ߊqw�M9��*T�i��kǩ�y �1�W�7�,�c�t�T��;/�<x ��O4�.o\r&v�H��h�\my�5��~�[�W�L�Oܻ�)����� �|8�9�|��jvI���؛)m7S7ӥ�Z�'�IF�x������e�z�C��>�}��`�}9I%���ì�����o�g�cX3�������ؼé����Ώ�F�[��i���2�+�0$�S�fR�z���B���C�#N���zPa}�l�>��ݽyAXW���QA�_�ek����b�ˆI���+E�T�s^�/��΂�[+��������l�T�kgD�Q�N�]���=a�g��8������fP+�6w6Yo�=�#:mт��<Y��C�'��d�#OR׵�Y�{���6�oe�4I���4|t,��O���*������](�]@��EѬDPCC��J���w�ZK�F�=N8%h�x�;�����o�&l��t���(d휢{��_�*3�~�֪HUPFC[�`���g��b�7�g�<P��u�ɡv����գ�Ϭ>'$�-�x��[`��f�U�����u�ހ���Hl�!t�!k��,8`ݎ����}���W1�N(�oM�&	�|���j��\�2��iw�2�F��B��@1�۝'I���v�;N<	}-�t;.N\�^��{cA���D	��\�8�\�?�K�]Eΐ��A����e���W7)k�s`cY�ޤTR��{;�($����v�Kb�:@.jd�Pwy���$�k9e���f6s8Sa��|���t�=O ���G ���_�$�gKO
1�.^ů��Xe8iHn�|��8��]o�Ն���)��@|����ξ�><gt�L?�S@^ʔY�aT`A니n<�P��*��>�E`̱�̵�	m�2t85	��x�^Zcz ��f)
L�1���*��m���Z��9�i��!n���H4�y.��� ����'�6YD��p�G�\�X�RNI/𵪯%�Nۿ`�-���� ����:V~U���x3w�m!r[��F���eRoL�����(t�JK�m�9�M�2�@�]������	b��5I���{a�y����!��c���j��cD�@�x�����k�;�{K:2��,�"_���D�J��y��AI
E��vቮŨ"uN�`�u>�oi�F�C�~���Ӕi�&�@C��ʏ��s�T�j#��s�dK�j�n+��e��#���zo�?�=��ⅴ=x��	Gᩳ_�f(|-���|?��׮�OJ�ԛ���Wљ�$ql(�I�x��&\u�#�|�i�'jsP�y����rydXO�`���'�_���'�_�3r7�x�䶢W�K����l�5�ȁo����6:&2.���K�������V�ho���Sc=�_��Iݐ�J��Gq�������˳#!N�#,����|�O�ؠ�88�h�z?'L��`���):K��G�n�c����n��";�U�
6��=�c�o0Xlf<//%��;�}���l�ʙ鿘��å��-;��̔�2;gl��776ZD�3@7��y�Z%���)�ӓ�3��		���5_��@U}�~�r۱f��V䱪o�pedzq�2k�t85�=ԓ���T�l'��6ϳo n}������,�s�,H��_�n�̊.�8���q��7�-����Ƙ�l�wta�5ke-�P��\3�U�$�" h#P�n'��`��x��aM��{55gX{�C���N�v�UM�.�Jt&������-���#�E�x�\��\��5�B�֞�s���7���H�Ū�X$4J��B��dU8#:Mi�а�7��5Oua�^�5%���o$��3�$�$�v��� ��$m2�Ag0[a=-܄�ڝӰ�~\�+ `~��^���_4п�+�<Elq��s�@�^�3^j�k�����`'F)0�à bNAŽ���!Ry�A���=�q%xsʁN.����J����n��~�����G&&�� �F�x,	^j��5���8��Vީ�>�I���`��\��-� e��'�҂?�u��20�t���\���t%q���Q�2�,0�+��!��=P��Xn��:��Uo�����m�3��u5����3�֔�ʩ+!�������+�ak{5����sѻ6�St��mo,b�Cy_@n��vc�3tc�b���z[����t������Gb4�P����k�W�����[���Rn:���$�S�kH�*�víb7� ��g�L��𢕺�w���g?�����7��(���6�U]���Q.m��1t��
Ы\0���4�?%;Rd*21w�ܘ�u��|tC�= �pb��Q���C� �c���ێ��f(\Z�~��O*�Mn���l�3v^�C��������L�+y�21��>�:�Ƭ�<ۗ/��pW��2�� .��G�}7�l��#���/@)F<����4��}�(q���Ϻ��"h�7�57j:o"���ᖭݐ[���5��u��c���c�t���,)�����K:��̕��K�L���G?�j�v
����"�V��P�6��Nc�Q��Ӓ�)�W��vp��L���W#���#b�I����Ine"�Xx��n�?M5=��p~�����ۏf���S&l�qqz%����t�=�?��ϑ=��ӟ�U۷�E�c�� +�d�������?,'�U�I(��	w:̞����x��IUZ7�I���j�"l�|��:��7�}�����U�i���d#����
u���08����xh�$,/����(�7H�m��08���m�)��Z�2�J�Q��>�.yL��R��`�7���m�~إ�W�v���ji�I�-����ED5Mg���Z�=?���^lټ���^�n�%��$[
�����t�t>w�ܽ�92�E�П�;�'uʃ{5t5��&��h>U��6ew�go�\�]��SA\8N�=�mL��S�`up�[qO�W��R��Sd��N�h<Rd�o�w�k"�b�y�8ʫ�\�VH�C��*��Y��a����/���v��u���L�#N�W�L|  Q쀱�����g�:E�^�w�|��&/W^("�Â�|��W;��b�ѳ�A��'��<2���q���}��C�`�ۥ���SOEx��M�"ɼ��_�i�� 0sm�ă`��sx�a�I���G6�^��=�to���}��wz��GG+^�!�����J����".A�Q���R�m�n�8�-�y�.\�  ��C�U�b�k�"��]��V���m-r]�H��B��[b�̐65�ae�%���]��=|���#+���%�.��,$���3�Z?��e�i���Q��xR�ȃK#�� �GMg���f8ki}RI�ɂ�Rӎ�˸�������Gk�c�8�OH1%:���A�{�W��rt�а44,�+�2@C)^;ӓ����l>��^�j�b§�
�:�O֓=m9�5y ��U����Q��
���#�`�f�����V+f�f�r��2.X�ΪCu�<��x�7�"b��������B'C�҂弯9�?��o�Ȳ�6Pv�	�p$j��2�˓���Um[�l߼+T7.d�N�^Y��~ 2�.��Sx?��hm�7���˞�6��e���["����F@�v'LA)�Q�xp����0~�T��5�ɯ1 �m�� �V},�~�o2��1�t���E��rI*��ێ�КgY�}y���Sr �.��@w����P�� )K �,�iCj�sG�򡸭"�(؜+�.�;չf��b�S�?��I�zJ��7��3M�Eak���Y"����wϓXQo|9hRM��[��gW���d�R A�](�}z`�V�F�r����ƫ%����{4��l�Ǹ����m����b���ۤ@�;���_)*�'�N0G�m>繥���C&lώ\E~�i�6B�#fXb�g�p�w;2�5�-�.�l��T ]^��狌����O��!�M@{�[A�qw��u�{nZd5al�L{v%��Č���
_�6��D���f��K�g�uGmx��˲��CW,��R�!����:��`�p?Q�����@���B�,3��w��U��*�n�^��cM�.G � HT�Ұ�5i����3���/�gPu�3�թ�Bf{&_���r�u|AÃ���SJ&��ĵ���|Q�:��k��X�4��Z�~݌����)�h���~����gP#��@��/y������)c�"��s
���p�4=�����ƞ���~W�����T�� q�%��5�m�ϭ�,T� ��=E��g��cq�=G�
Ё��Mk-.�,�&��ѭm�Tl�Ӫ��ye�6J.�� �?Nu�WzXf�N���=��������o�_J�l�W�;Y���ii�-��]���c ��/��GmJ��j��"�!�5X����T�`bF�d��A�R �p�m�b��牋����w:D������곘�_�k�����;� �����7��.����M� RF��g����i�V=�rV
�VbY5��K�:8)B���/��Mw0��o��kiAx^��B�@{������/����T<z~���s��H/��1{'������vs_N> +�=~�v��f>m�w���>�֏���g�{����M�����Z����M!������y��gK����q�Z53��q��Ǝ�����:Ig�e^)��8ڱ����=T���f� b����;�L2�������ћ(�87�{6���&������&��<N��'< �1�����`�[[U�ɸ���YC����is�ZC+�B��~����d���x�����r��A�ϙ;��ȧ�A�me����y�oƳ��2B���RT���>%O:_l�6�;k1;M�Aڈ�t�9�赉��Y�3�VV�=u�&kT��W���5&ژ�^����M��TZ-'�Z����?k 541ԍ��U��*d)Y�)�zj�/V\c!	��s>� x�40�Va'���v+���C¯����c-&@�#Վ_<	1���&I%|����z>�z��hG-<�ѿܙ+�VD�bف/T�U�;�|E���&�xoޥ9��Zh��q�UM��Z����.qm�u8���=*����NY�L451Sc�k|�tLam��EeŢ�w(@B�S�z���ݘ���<�н�6�e���=�E��.r��)7cE�*��5��u��ށ��*+�l�{ߦ$������$Q�akE�J+կ�������+�+$O��N������˹�^
�����#pk�������?�s�;���G�I`�6� ��'2�!�׺�[n������taH>�����ه I�% ��!��5/榕��l�t0<�����Y�@�!��8�Q���Y�>l\#�2r�;#��_�\�y��F�|��?�T(�|�Jc(|"ek(�������
�&."���,dq��_�Z��������e���Σ�����d�,�&ɀ�^�F/�Aփ����j�w��$[��5���h�k�Q�5��#����>R��Y���"����D�ʼ�{�z�`��䧸��S�WB���;>3s�k����_qmT��uF��� ������4�7J�S������������{����u���W�v�q�XC0��m�1��ǵX~�3|�����폥/�ʹ���1��!CV�5�B����·UA���t���ND⃶��fR{��/�ie�/���ʰ�q"/����hKn�����v}�Ư��U|�Л3]� ط*w�5Kf{?;��@0H\Kr~�A��N��"9+�-������ߢ8������޿���O��At|pDD��f���'���.��.@r��O:��_�堳2)g�9�,�v|#�zl�2h.`�5���S����D���od�8����K~h�۟5�}j��J_ �������5�Nf��\�����_Cg��e�����N�2i?�_�_�]��Lm��Im�I0�;�f�-z����ZW[ID�(dd�'�r��� $g�߅tˇ��[���uЉB9;�^k7�
��Vi��\{�����{都�.|43~��Q��"HwA��F�*(H�ދ�( m��! -�^�ނ�@�QZ��=%����?�_w�u��Yk<9���.�~�~ߜsR0{��>]�O���*���9'W�E�U���6#�#�E �Z��y�tj��IEN�G�~�s[��?�f��Ku���{�t��o�A�"��,��D�B'y��rƉ�ݾ�ވ�j�g�U���r����#�A�����_�R�i�Fq�s����Ŭ�(�\���!r�O��ǚRW�98Lk��� ��KL�AP֔�y�}��a��\�~yQ�3t��-)�Ϟ���_42o�'��-B8u���8g�@Z��D�N~�*���qЃ�Frt�A9��R�n+�#d�����oE쓧Y8ߪ����8Fg�,��<��Skd��p�WS��r�����k�f~�	�����{+��&'�����h3��.���Hea�p_$�B!♂���rY�vS},�QD��!��i,T��:H=�nչF��U��6WG�~��H�ͱ��Vϼ"�9��YcN?���:���x �l%Dy[g��F����r�g?0#�>�ꭔ�'��1f�ӛ���j+��=̡��da˫���{�Ǉw�'!��D��5�)��Q`dY}�?��Qn���C�"���  �1��8 y��i����۸`c:�s���a���K2�:(5]����יQ�5|V�oKa|��K	u@\YZ�M���G�)�����|H�m�T_OW�mݿ�+5�Jҋ�sx�r�!�ʟ�R��u����v׼b4�5��tF��c�5F��)H�8ʪ�V�̖�U6n(���Ӹ�-ڧ~�? kU�i���b�"�2�_v��n���?��'��ʟ+���2Dq��o;�G{��)ɮ���Z���G��&Wȭ�#Pfl��*j��xO�b���G,�
Jl�)��Y6����;Q�W)�^=ao�I|i	�D���ҩX,��E!9n��g1��l�]`d�zPV��Ā��*��F���k��`A� .��%���zf>I��)V�5�ȟd7�n 
%k-��BI�#�B��fx"1Ů$J����@�c���B�mwM�	x,�qq�m��u0;��˥�N��9�2͐��YͳTV|��T��,z�\d*v y��wg�{E����׈U�D�OW����
4�/�o���@V��$�{�*FmY�r�Uv���pZJ;���#����}�jH+��U�����:.(�I�䷪o1'�3hUt$F�۷�I�3Tؖ5B�K���/b�]�g�/�B��~�|WF��)��;�`e��y�%���0iw�IĊ��� �͙���ѣ�X]�uM�IS~&�Gtw�g�N�	�Ո<vK>IL�pn��>8�z�։���"�o�UYU��S	��o��)�L�Y�W���t/}�>�=C�@`}@�� ��dv��t��s��_1+W�Re3J�>_F��8��4Q
���o	�F�O-��FFc�zF1�ԗ��x�u�݉	�SԽg��	�jE�S,�?��t	=�򕉚��fz�ߌ+7��߻ᗃ,�,hyfT��Y���,p�r*��3�]g: ���G&NIBn1�VÞp�������4��$~���rU���G-�29�{�\3�8�J5�k�a{)̊�r�^.j�.x����J���8F�tX�"���� ��$u����$�� ���I��x�+W�Ӕ���.���� z>��ܾ���<���#�
\+7'>����Ox�w�]�߼����~�B�����f����8)�S��r#3�V<{�۱R��t�KÊ�����YNn�g={��9�KUB�c���{�G�G�Y�H���ouM�� Y(�^Vڃ+�q���oZo�c��=�Q�.�jԛd)���H#$��	r�#�l�$�"{\��5*2dX�����U������|��?{�f��
`'�lN�9�r$�0�m��҅�$;�r��=��0ҺY�aeuLo��&Y1!n��)�s�W��tS��>!��	.&>~v�1��+�?P�K�Q��{�얺�u��SV3ho틍y�#-a��>��*�V���@vm��L/M+��@�Sr�Kesk307;F�W�>��������Bkc�}�����E]ԒӸ�Cg,3����v��1�q�����3+~�*�Q�{Z�]�~Yh�����w�!��&���֬�(@ղ�'VzJ�e�K@H��@_���Oֺ�Oo�e�I��avT�����(����_��WE�,�)���ԟ�v���?y]]���v�[=���7�Z����o��U�,�+Z����;~��~pk�peeWNˤ�tk�.�����8�+q�3po�����.{�J�a�v� �� �#���tWxzv�54�B98���m�"U�W\C�@��^��1/CW�i5c����S1�}����Y�	�J ���.ӿ*2��:�����s�q�х<��)�l73�,pK�p�+���c��R]�{���3���w��K[��T���k��KՊP�LMWsC=;���s}���i�tl� �&7����q�c�g����Q�l�y�g_�K�^-�������`������m��wW�k�r��e/�U7ơ|���O��S�o/w6٦���|�Q�n�飧�*��T��aq>S�,�";J�k���-�ǎp�_c ����ےd������F��"w�s��<!�!���8���W_��Ԍ�xδ6V��E��=o27s;��V��B�A����G���U��*:HSz10�H3@�nlՆa�	h]ɍ!�mک��&kooKY�|8VF`;�*��H�������%��`p�'Ǘoh��^Ff�&����`�{���[;%X�Gܒ�.:_2�^��2��u�9H`��'	�<�C]ɽw-Q��i�� �k�����+g[�B�S���Wf��	��+�8H܍I��.⣳�ՉE.6�O��;/ϕ����Z<|�{���ڢD[�/�y�>�c:ut���RǊ�����j=	g���0��X[$/�O�j ����������
�����b�$7b��4�2��ţ�X��b�v�d�z��'�j�H���T+�@�o�7��"r��H���ys��$6g���eO5S�/�a�X2ʗ�I��dU��b�,��x�b�hF�Y֞�"�K/K|	�5�K	*vb�K؈�����^����o��lx˄�_-N �}�q�	���0I3�9�S|w�n��<��뜅邻 ��e%M���jG�ṡ�[O} ��Xg������m
���(ɝ;,?`�-B򐔧�xT�� U^$oa(N@B�_���b��zCA��^%b��-������w��J��K�-� �TV
�6jƃ��)�Ȱ��fc+�Aޱ��q\��_�.�kg*$2���ܖ:q롷�(?���󀊖��E�d^��=���(��F�׺������.X���l�Z�=�t��"�5L���{�oS��+�o@��v8��X�2��DUZ��K��x����K+��j����b<)~���<-�'^f���s˝���G8H�ɟ�����֤`���`�Z���|�;�^�hF�۩k��[N�	�\Tϧ�|���yϏ��gGqdl�\���bm!�Vda� ���O�j�8@�֫����=�*�u�R̍@��y`�&�����p�*���k��`w���p�jk�>�"Sġf�@7>*[̿��a^Ü��޽Ԟ���^�o`P�t�ʊ����W�+<���1_��}�7Fy�J#� ���Ү֝�O�;�I���,�[[�؝&��ƛ���̷;�Ag��D��admQ7����&%���x�8��qL�v7Bq�n�#�H���c{�uA��0�� $"��v	�fI�[�T9�6^�:�~����~F �3��Kx�ȈDh@�)"���<���SMd}%N�kn>X����g 5}�+W����Rܜ�����v}}�����֕Sl9 	&K��O���C$�+��k�_�dv��ZP�V��}�n��Ħr���P���:�sR'�g��i= �"���J��{9�0��_�,����^qu���-��B�y��W�UX��S��� 
��6�}�~Q�TЍ�5sn0Y��07D�O�e��P��'�v�&�H��.��f���7�3x���<m�n�`�1_KE�Y@�����$�T3�mGB7����/{��u}�pMD��)����+�Z����x����!�(�:��@���Op�¿� T%ɼ��[_M��� �
LT�l]#.��6��6bv�R=�?X�|�0r��+�� b��������zS�(�k�%5H�ۡ�i�����2�C�KK�+l`�IRTT�0gt�����ػ~���ot4A���pQ��?�@h�Pcִ��[����t�b��������3cAlxF��i�l��#��B/fB��J����;H�-..FAij�ɐ�@��е�$G���-z��tj�E`n�]^x�b@�)\PPi�Ę$��x㨈z]�
!A��{�[mv|n/�3�rm&��u�����C�N䕑�g6�U��n��Cg�6ϕK���j��ޢm���o�3�-Sɡ���9Bl+�K9���2��¨�h^���*�5��V������n��0i3]
��=M'�����'!͟�)ߒ�J�j	�
o�:6���>R�� !Įnq>`{9H!Դj|o]M_�>�m-��N#YJpr~ZoD���zO1�s�g��_+=���^���qvވ�&���)�}�ͫQtp������n(V:�r#�k�_;��g�������T��S	�v�����C�4pa^/YUU����!�SnÕ���m�h��+={��+��H�C�L�3q��p7R�btX��pKt�y ��D#P�_�9��e����ˠ[��w��+�/҇5�&t��Y�농g�O�UK�Totуޘx�v�1��m��|���*{;�����RN�u5��S�LU±o���9E�Y���V��٘2,j�����1��!�1y|V!��I����z�|U[�G��7�͜;�g� Ă(���m~��t���ݾ�<ohlh4�w�ٕ	�5F�'�>�䊬�oo�3��U��ʣf��:��|"�rdׯ�	]cN�nq����3�UܲE܁q$s��׼�� �G��t���$�;�lT�1֯rZ��3�"T��S���z˙�n�7���~��)P��F*�������z!��#��C��G�z"Q�a���R]�m��:��-+#I��Kń�g�Y|9��Α>M/�\�\XR��� ��s��R�&���w􆉣��3��Q�2��@O#��-���I�-�ܫ�4�֔fsȧ�'��ax)�0`*D��x����^b��7B,�g��l��D/t��Vk~d���E�3����7X�-NUpj�o4��G�2
' OK��{��1��5�������P�}���\o�zn�z#��/JA~��a��kIto�+虚K}��Qg��݆���9��u��7�֗A��;7��7h��s�܊4azl+�Ѻ�/���f"�f�y4��hPE�@+:\Z���7k�!0X���F��$��b._U_���Y�p�JHk�����0�%ZH��Y���r1Q>�3���@�:��3Hf�.�NvHc��/O�D�8EÁv���ߗ!A�������#c����0�!�S�H�@�
�2�䢇���bE��0&s�x���_�l۽�3}���﹑7�#�c}��s������wC"�J������z��[-���A�g�`p�`��2L�>��������,�p!H�/��"�;+��-�$6`4���wD��jj��1�+�J�m]��iy^�QJ��}�c�9:�,��kjC,�2��Gn����V%���i�Í8�N�׍�;�V�B̜��T��=}:��RbފdT}������Ky2���P~� �F}b�zI⢝��b����"xiW��FmU A�����\�W�J_���-De�ˬ�+�u_���q�T8G'��M����J�։ !�K�!���FE�+���my����1�Ӆ*w!��i���,H�	�>���z���u�^�zc�Y�ż���g���n�us��ZGsWY�	m�Qm�n�hTp�a��o���wCu�Qs=y����@k!(XE9��~�ss�PHz\&/�{���m���C]T�{V	�\R-sƱ=P�'��w`5���|���y�_���B��M˛p�0��l�a��V����8�=�����M��n�De�@�Ǐ`󆧌��Oon�{�s Ȕ�r����/r��P�WCȌ����4������Ό�������QG�_��NȘ�8a�'{�v/��%P���F۞��+�0��i�}U�0��z��x�����mC�� �ăN�q8K����v����1˽���D����|��̈́K�P���w�'�% S�w��CVJݯ������7���/�+y&�����k�y�X_Uܢ?@s_� t��]�_f\u�Զ�Si��L/����q'�5>���D鍻y����@/˥1��'Ry�|9��r�α���264v�48J�ɽ�g���o�*���vns;�2�:��e���- ���x�wo�a�Ҍ�ǃ_�H��j���Xy]��o]�W�>w���z��}�07竐�6�6��]��.b8�nl��|�m�:$��6-����^�o�N��ꘌ��_!�8BL�w~��k�el���N�v����I�yE3��7��n#7�{t-�z|�ɯ��Ef����CU~�7ꣃ��� w�H��"�^l=ȇIf��Աl]#*?�t�p�5��lҘ�#�8�ߴ�9�Խ����=��� ��'�1/#�{�q=������j�K��+vt�;��À���}׼�ja�Ѐ$s؆�|��=��Ώ�_��6��sx&��Eu�ӯ�/8j^��]/�ڸUW���s�j�vz}r�6L_���q7$�-<Ȝ��s��xQ�yH3�Xܘ�ĵ*Q�y;���6����6�/�B8�1z�"Wc�YQ�k�4q����H��w@<��f������1�1�����c9�}�
��Y&�F�@�y�ck",+!G��.�&C�÷lw���K<��x�l������;�贈�V� ���-\���k�~:䎝䁈%G�P���,�N�k����ޞ�.�0���%�undf��dn]��a�Y�g`���܋���>� mb��8cl�A��~������;�o�/�&�jx�6�]�] Uj:�~�]6IL�"��9魕��M�J�Qq�.�n�*R��e�|�3u�Vi�s����K�Y!�m�D ��[u��$��7����'�.o���F��*�ް����Sޡ����	���1�����N� �W�=/8���إ$���%�
�G��4Qf�A�Q�՛B���E7�r[<���fm�.?��������{�|���IN{IgU�f��%_�d�s�jG�w�0��������S�+OA�O9q��q��G�Sϴ1�4On��7���M�j�� ��x�TJ�[���&�<G��~���
d4�3cX��� �Ȇ�z<�LUL�&b�������W�hX䖔!6��{�{T�~mÆ��>j�0����r�_�"�(���I�fO�2 �z_!@NW�}��q�_>������~��O3����y�ȷ>i���6��e�9�V��)����
n�*�h ��̍��&G��>Fa!S��/~4@��n��9G[>��/�xz���ӹa����?�1�Z�B���BzC̤,��������S@R��&ō>��]N�
��g��ٚ�j��F�tGo��*�f���j�xׄ#0+��ж�m��zȤ�V�2R��k��=X���?��X� �E�/^�{^�iqQVD�d{�?��n�����cS�U`[����RĤ�S ��TR��8�����'$(��X�"Xok���u}�D�����\�,bp��h�A����@hй�����0������]����h����Y�X�_����Ӣ@�X�rX$�x���%��c�XԓUOeL,G��-cօ��Z���(�	3Z����~�����v����V�3���@���0$(�X��_\�Z���}T��﷫��G: �a^��$���F~B�g��m`Dٌ�N[w�<?_������m"�\�q	׀>�g��z��O��3�'���
��s+�Iw����QT��P@c�� �_�}���@�h�g����|"}}|��i��0t���" ,DH�vC�ר���k���:��Æ=7ȮPle&�L�*ف
u�����RX݀��z�����β��>;�@�)�:�l��XK�������N�:gC��`1�5����
u�;c�#� �1}9�U���~h׫�6���Z��������f<����c�[g�i�0$�-,��ĵ�Ny���zR'�4�Fݎ��� Z
��\�G�$!Ɛ������-�p�� ��J1&Zz�/Vzz���ֿ�X���]T�-���/����l��sk,��D^����x�ǟ�3�K�^��N�;�x-���os�sq������g��-d���W�y�1�rY��e��	L����fW�&���!{��w7[�\QU6��]�@�^�s����ƞd#��R> 㤷Q�e�����
!�(����	�)}2g���!Q#��C�c����X\E���Q�h�������5��kR1cvc�e�� ��C͹Ț*��N�-AX�I)�cs��*�ƈ��P�Y⑪�Y�#��+��tga�j�[z�2������;oA�DM�Jc��4y���V��cJ�O�C��[ ^]���U�;���8�6GX��;�&����$�H�Ϳ�y#��b����t�e�b"�탠�P��bn�ǌ�x��X�7��yW�)��=��=�˭ixP�-�T��L�閧i�G�d���6I�67�� �o�nxb�t�����I�6FY���l,�=4';n,�`��w��_�U�+%�Bum�m�o����=�#�b��노�"j��\�)�'t����k��O�&=�f���@tq�YB_���w�K?8{�v*cF���gq�!j��eg��<���D�\�����3	|ԏ,}���r������p������k'K'Y�5�\G4�KՃFF�d�"!J�j5n_���V�]FS�����l�����>����hw�Ul����k_�Ұ!����w����)v�G�v�� ��HN����2��:�8NK\1�gU&ħ���I��L珙�#|�~`#��򄇮�θ���9$PTB���H���eU��E�jם���[ë���1W�_��^}�m�D�._H&���)�I]���݊M�`��K�J�+#d�W�^������@�ę�lժ-�u�~�iy�nk�w���W�'V�OGlW���[�5`���d牶jhO������XD�� ����;��rQÿw����MN�\����*�K�A ؽ������yF�yɮ�0�	11-��?����!�W_�����m�f�cϘ�y�r��?d��[���7O 
�C��`�_i��Ǝ:fo�*ҝմĺ^��cc�=b��J�����!��e)�t�c8w*Q��d2�HT #2i��9�zȫ̲Z�'#%C��*���ٮ��8[X�*�T�_�p!�2��^�I������ٟ���>h�����������ܵ�MJ�~���Y�㐴��Rl���H�4A*��t}a�����9�Uy��]��e��o��%�U/����vi���5����i����Y2�'��C-�S	T����\�)�A��tS}��ݱ�;�`uu���li�Ets�]��x@�j^9o�.o�D��ƪ>��,�|��,ż��'�m��&g�#g���XL���R���S��� �:��)�a���o�@�����j���6�4�R���w�;�AJ�4�@��&��6�98��E	��4��f��H�ʉ�PI��R$���W\5�ζ�	�؍U��z}D�K��ꡆX�-6s4g�b�mb���.Q�6ѷd:̵��dT��O��xɼ�,6l�-��͏�p �vM�F��a�cņ�0�����s�`�E6�ա�\�X�/�zyM��j��Ʈ�TE��ϙ��|y��+�ٮ�����1�N��F�}2�n&B�"��t��D���l1ks�Ғ�T��5
6���C$�1*0b�3���np����̋X͋{"�(��<��P�� ��e�����Uk����I�,�t35^�_��U(Y����/]ƃ�FË�y����fG�=*��8��Ƴ0���5T4�y���� l�*���X�X�]Qܽ�:,,e՟Ӓ��M7[w�	!�a(���/o����\�Y�u�x��J�i<T{aۗD`��3�DW������r�=ҕR��[\��CSyR�ƺ¬�t��+�}�Xgn��䎱�Θ����0��hv�Hh��[��ޅ�����Ǭ�;�n��Z�����R�-�М�)o{��'�)���kLJ��%]!Zx-߼�Rl�#b�#�:��}���~��Cp܆ +�д��e���fѣF�P�Pj2�^�c1a7;f�&�ی��.�F�i�yvʰS����G:s��Ꭲ�����t~���6V�M���B�Fkqp���C�����B^���E
���zwF�z�}d1�L�.�(�y��x����~�5m�?oT.95��!�D[n�"]#��.7�@"_��}�f�3n��q����X��C\�S��!�@S^G�p��@�#(��z��[�5zn�;�]ݓ��g3���Xm�9����06�~�2e�dAiX��1�w��r�Ň߳����d��<�����7ǨwW��kC�H��U�4/��ʒ^U�8�zw�:��࢛G��vI�j|߷R�x�Q��{��#̽�!.W;D��RgR*���z�e?�b8o4���5��</\�����m��k��a>9�lpw!�z�SP�Fa�n���j�a[��� 1���Qo l�˩�4V7��	P,��V�L��0Ow�f����xԏ�_��oPN��(C��bO�/�	4g6|��Qu�u�¡{l���d���CA�MFv�?�[R�<]h��H��_�\���n�8���:/%P��X[gZ�34=S�c�Q�Va�fr2w�}R�%qaOD�ce��a�n�?��`u=-˷5Rc�x�dو�L����w�	��K�����,w*=�.6��ۮ�Uo�&xb��Ʈ[QU�iO�O߬ߏ��s(f�j�mh/86(˼m9�.o����t�=��C8e��ZԱ¶�B�ٻ���eݹk�:r�wP���쀐}U]�q=��2�� �ePUB�=�,T;#���'Kץ��*ܟ����;쟕�X�>|�-���f�k�|�Y<��|*�|;�u��E�����_'��Y+g�ެ������,>�a�ݺ�{���;�y9rAw��Qd^o���n��ey>Z����h 3v���^$���{�?��W�Vǖmk�9�ʪ������L+��E��d�	�^k+��OV���d�>�~�ˣ���v���y�p(zV�6`�m������O����{�b���BZ�����T�eX�m�+9��]0��J�+�t����Pf��XY6G(u��09�+d+9Y�b�ꄍ�Yloj��a�3���:��������=��d��r�����	���%�:p#/�G��7k��U���S��ݑUO)voB���FJ��it����w�{��{�a�C���~���1����\1��p챫!��g��Q�(9��ȅ���ʬ���v��d������1k���c"�s�±���e�N���կݰq5W�-  ��QNU��jrvB��X���-���������U\�N����bY�e���}���5,��tGxu�Y��Tx�R���S� C�� -h�})����'���~��q���'��q����'ݐF޴{�?�܏�?N�8��䏓���\��B߰���ۍ�^������?�~�8�q����я�G?�~�8�q����я�G?�~����'���Kb��wuU0�����tR�׶+�O�Ҝ�t����'-/�oӇ�'䜫°Hޯ߼�uH�Th��~��%��OWj޲�_�RkP8]� t���W�YUħ+��v����z,��w����[ۨ5�_�~���߻|�����
����5��9���C�?�gK��c+���D;Hl�3����cW�;�[c�E�.<���w��+���.�#Q��P~\ $J����W�=T����D���X��Lm�����?%�1@׼`�9al��Ο[�o
.WP���i.��o�W��R�7ܟ?���25=@�q�',:}2be�V�7�}�p[�T���'Ta�B5w�C�z�tA�o��������ރ�,�'h���E�^�
�>���w����4��ݮ�A��2޷!.**J�������P�F������!�ŕ��r-�2&E�@�qG�{N�w_3�u�J� Xrξd�u3�������t?vѶ�nl�ݿY�٤ؿ����X 3���b)���1]t\��)UƓ}�
�A��p�j���OA�u��ut�����ӄE~7�2v�����oǝ��2l�j�����
�϶���X���4� i�?�]H.yc����Rkʻ���VAl2A�%f����GI'c�<�Pj��nh��G�[E4�"EUuuu��ak�������W���}?{�:;ĕW�P�<�!�"4"Gb߉��)&���s��%<�mM�87���($婉��r'$���L�Mvy�:�w����S!uMfߓ]�����*�M9��=�]
�ː���+㱌��ꎷ�^4��d��J�f�
��+L�tH-��t�20�^���8'At�hk;����q������	�a 	�<j׃���y�o_�%(~&Vk�U�kY����@@�\*	Z::�gXA�֐��z�x��S�����!�V�[O-�Pe�>�9��f�xxx�
������K	��� ���b�)F5_%�o��뉚���:}����5�wzy�i�@�;�������˷wv]W�o]�i7��W�p�:J"�o�Rr�� 3�333P�e�QLy�i�#�5&���8[���v�$t���:�P6��e�/�W��i�+VGԨ4KT�cg!��r�n�	�M�B�{�vή�����H�ґ���X@��(d�����k�uThzH2���L�����]G;nb����:�/�TT� ������\c�cs�(U3���Z5>�+PJ��W� ����a����E�n��r�Q3�e�O)D�\g~~~�<����4�ɡ+$ O��;@Ss�
\��@���~�vUA�]5���7� ��\.��B7��@��<��/{U�Q�~Z"�H3������_ ����s��tv�`��]|���!��?�/W <>svH�fr��xG���:} �j���DӜ�۾��]�j��ffJs�W�ڿ�[5~G�淀�-���PSSs}9�aߡh���ȉY ���D���PSB�\����0����g���a0�q�D��)��./(Xۄ��˚�S#@��8���Y�ͥo� ��i��%�#SG�����02�h<�0 #����q����Xg�DONø���x���%����]�=��!p �>�̖�p�c]7\*.��ߟ���9k4��9�'�XMHF��CT�@N2���@Q\���i�@��@<��~��;6P���Ls�R���%ԣ��ɭ�pӵ�W�A�6 p���B��09�M���Oi�>hb��-U%�EyI��>�f��!��ζT�3��9�c
j}�Ga�V��!�f6�x$=Х��㱫�{w��	�TKO���C&��QB�U��~Ԧ�&%-�����Cb�u۴���IN����$���É!O������V	93KK,�L���O�Q{��W4�
S�{Z�L �� x�WdA��y�WZ`oz�9���A�?x 'X[[[�|O@/<4��z�+M����g�����Th*fȲ18��P�v��A҄��my����n��z������	Oy`��e�N��in�x�wK#jiU"|ͥ����˘�L���Rz,�2�<Oʞ@r��/ W�`[�[�E~0��!/�H�F�("�9)������p�Ҡ�#�b�Ă�oY{�Z�0�}W--�����F�8|��3���c�T5A�Z�]�J،7U��}���0|���$��K�
_n��I�ﶴ�S���+�"�!11`�zW]U���_v�Z�u<�<X`.&x����cN[�s}��<
�4ʶ@�@��`N[`���չ���av���"hN䔑�@�_�ψb��`we���}�U �&|�Y�Fu�W���F�E|�=��^��ȗ�y�@8����pD>�][d�p� v��c��n�#Ǥly��`�lQ{[���
��#���7L��,-�"T�Q�g����Z� ՗�ke���&1��[@mX�<���%�6�$`8�ځ?���#�����d��@�Z��#�}_6Ix
c�%����,""��{�z����j>��- _<&:�8���Q��aa�!�@>���[QV�1�i�3m�EcژP�,3�3�x#cc��Z�u-K���$7P����'����u��m8����aB���f�2b�X���c���c��J�K��[�a#vz�0��ɖ��	���67�Z�sI X�U�A��7B+ġ0�*�2�݉�86m�Y0���Cb��|�Ɋ�.Yba��i���wIu�h#	���4ʹ�`�4�ʰ�P�/����0=�#1� @��n�E�>�e)�D8�\��)�Y�xR��Bf[FO��8S_�&����r�(EV����-�� ����#u�ڄ�S5O�f=Z׈F5�����K��7���H����ճqp�c!T�j�^N�uX)9y芐F�dM-�r.l�Na��5��iJ�4_���0&(�m:�u
5�2�����IE3��f�2�bꞽi4��zD�꾆��iH�	=��c}�
�I�^�4�ޛ.w�!�|���BzG�8���g��D�6+ ڹH��^�Jo����1�)/h�؜<q[���P4dL������n5N4�����
Cm�slQH�H {����v�kceilE/A� �������j�F0��G;��(3��j�a�8�ٙ���r�X��kC/Vk*\�AՈ�	=��G����4O"a�rv�&T?qvޚ�Sߎ�:�1,ú:����>�pqw߽� Ʈ��f]�yI�)%$FĆ���a�L533s���̯��$���@�E|c+
F0�6&�$Z]aUCID��Mڧ݇}�P�|���X��������U�Z.h���A�a���p�s)���C� ���Eh���u�$!"��QR���"
��аk�/� �!�/�v��j^"�F���JX�q��i�z]�*$_zHz&	�	��&&�H����*r#3+�R
���;>��7�c��q�C<u���˦�W�"+���t'��tͯ�3�Q+��Ht� �����+�2��,%�*�J��Vbh�:���=�bʶ����j�WZ�)f��<�e0X�v��?M�0��@�L�Л�U���(8�NT(�Z���T�e�u�����~�L��_�Q�/V~��� �gkjk��A��&��*�c8�th�J����k��<i���73$�\[N���qqo���kZ&y}�!�"��A��t�- ����/fh[o5��9��_Eb�	���X��N�!mw����E᠋x��;��Eߜ�O�iha1���W��}Ti�I�1�m���j�J���bB� �z5�huw`ѶϘ��V0��E�Uھ�W����2	�s�@l��Ʈ�v����N�=��Za���+P�a�3Qê����~&O8��S�I�Pl���4�8BǶs9�
��:�f��b�馪� ҆ݑ ��	}zBX�����~�����5�]�;؀E^V�Ÿ�,}�%�t%GC?'���BZ���n�^DD$;����H��`^�\c���ڃ��gˢ� �O}N`��.H7�Q���Pl�6@������,�F�q���dES>����⌚N��0t����oP�hL�{(g�����L�Gmg�"b�v���WWW���`%�o��q�×�GD,�!��B�<�!�k��O��}}r9yy6$h�Hj���>ͭR�_1��x�e�i�����%XM�{�5�gz�-��W�zIV�ѓߠ 	*Ӕ�VD�o�^�Q	ڏ���(��54|����Z������@�^����F�����v3�,Q���=
�.Z��={V6¶
�_�$�cF(|߷���t����t�vQ�b w\���istPp�՝��=999�n��x���
�nA�������u�H����К��O+Դ-��C���n�AY^�8�״	x����!_\_ ' C�m�}�g_ҹ}�z��d!U���Zn���^��[˕���!�Or(�
���b0b��k4d�Β�>X*"n#ו�V�7
1��YA?�ѐ�-lp<�AZek=7��ߖ,�Q��(�"1٠��Y�<v)�/5���� �͡h����{_������^�,m�9�tb����[)��[�"�R������Ό ����~��nn�@>��� �	�cCb�f���!x3=����1�����p[��:��B��>m%%o]ϊ`�� ��X�=R�h�������� �:X���$�E*J .�.��x/�Zu�t�#!&�|�Pt�aoЖ�\8�]�@�>@9�,�[��8���sh5��V��tr�JZ�I<܍t�RS�C!+%��Z�B�a����_NҺM_{�q'5�+���(	"OL�$�>M� �M� %��A��PfD��2�����(����sK
ͳ��\�QS���G۟}�S
��ǋ�􈣥G]LBB5?f�PV���p[!�U�F�֢_��q|m�!��$m�A&p��iN�m{���0СZv�}���5���2�XLF��ZB�ދ���nF��M��?$���M�Du�Š�����P~�����Id�fmT~�2F[P\��7w���@�%��E������ȉR����u)-�@�����_h�7$9+�0A������`��x�A����`�bQhW+��8<�;&TU\yuB:��b�t�f�uz��N��Ih˰$�h�f�Ä�Ā��g������L�C������;�U
�����ܭ�H���1�9��}�EX�EK�%�/ ���ښ�o�Z*��ּ �2B�g��(�� 5��hn[��)��AVD�|�Am�9`a�]�4G@�U8��cͥ���	���D����i\����W+^��*ⶀ�dorX�AK�:}��v�f�*�ס8@Y;DOu�f �2M�D$�E���R���@_���V��[( �2�1��ͩ8t2�*��3��CGN�qb�V@��K~�*qe@����HuF��XNP3Ρ����((X+�L��` <���tP�@�P �4�62��q�)'4I$R�P���}��䙲*���RrmIV�{�FB�-W�W�?�o\oV�C��
_�K��Ÿ���o���x+E��r�7�*x�'Atc��s(M�4�����n{]7���5UKg(|t�Q�_�q��t�g�+���ڈC�l�W;�e�}G^�ԼB6-������݆	\#�JcQ� ,b�A�zL2g�1ڨ5�O(���$Z�M�f�}�
�6Z+v�/I1h�\ޭ d���@?����˦�«߀6����=��/�c/ɐS��t��N/�A7�6Kbo�voĮ`���6�JKK��X�^HHIm�%"�/��@vz�{�!�xy?΢S^��Fݕ�U��pq`�@��k�ɏ�K+�qژd���8h�(?��n���R�5O�VA�_V���%M�'��u�����k���9\��r�r��c��=z�h���
 �ZPc'DW Ovz
p��'�����D ��и5��q�_�i��9�F�bP$���ï#@��o ��2e'YMO�������#�)�
�s�h���*I�|0\LMt�h_($)�����n;�.�����?V`��j(�΃�;%N� i%������� ҭ�mG�����ǽk����H���nAU՞!�2�]�-ԴDR��Faa�7<0o�þu�x��Y�R����[�c�A�ʼ��H8h��T�?����˩�0n�N�1��j�(!�ۉ���C�=E9�>��^������S�&T�A�7c���v�I��J����hh��G5
'jk���P�ǕcT2�
�#�t��Z{,��5��nՅ 9^��St�����;�ɫ�?�����jS�� lhՈH�( ˶l�XD�.(�e�n}�("�0��*�P���(2D$�a�BD���s��<���W%7��s��|�x�s�vOll�B�j�{Fz':��?��<��d�;�n���444b�+�%����S�4��I������#��K��b� 	���ÿ�1V��ד����fRՃrL�z�#͡�Z����?�o�M��!���%��q���!;���5���[+�kF���H�讋�6k�� �ʡ�Y��<����Zz�^=��	n4���2����S/�}������ݙ<�@����O��.�C��8@���'�b�) �Z�L����㣦2kz���JR�*u����c��7�V�d�d�$�*\I�P�Ɲ;���5Zx�~_���w58�¬1R5�*�Aro ���bV�*���Z�K1
p\o��U�g�����X y·zRC �Z�П;0��%onV���V������'TH'	� ܲsR'�i�8O��¾M���P����<���6~&���j���#GV����r�V�\@r670��X3��U�{{F��]'�q�npE&%W9���Em���G�n.6@2ʉ߁QTOp%��A�HQ'�3�º/b&yi��F1Z�8�c���}O��l羾��Й$����\>����B�J{�y��م�$����>m�9p�߷5Ҁ����#߷Ot�2J�J­�֨��"B��B�`���_�%|#��d��r��z�w����њ�α��X9ڴ�{`�J�vrF�w��S�]C̽�+�8���[$���߹�I�L��I����>{oi�iIf,J񕖝�m��]�ï�YkH�Y��N^ ���d� )/|�/�R�dX��St,Z�`�ĭ-i}�@���N{r��SʟlXЖn�����,� d8�/�������+���2WB�G���ca�W���U���lv��T\�� �	0U$����F��1{NG$��s���4H�3\m���XQ�v�n����$��~�2ؿ��<���`!g%�SH6DtY'�7sETɅ ?%��1ɴ	���F�1��������?|�E�䐇Ė>���b�j�m�qP�+�+	�&������qݑi��,�ͽ���
P'��Ha��w�f�;;��<<�� $�Yӵ �f�3ݳ��.{��o��E鶧�Ѝ�+�����9&�p����~�,�ـY�G֬��qf)��xtZ}>2-a���@�f+G ��͜�\b ُb��������+:F��j�p.���� 6�Nn�솵��O^��e�6�����J�
�H���w� �RsK hY�����>,e!���f��;��Vlc�:�n=�
R]�!�[H��N�Ž���J�қ�-j�$<�:����VO���S�;����E{ƒ ��Y�F�ϥY��L�z{�!�F ��S�o���=��B�!������E�����б�F�r|F�pV}�gs/d+ʊl���C��M�ʳ
	�,��@�Y�Vг-P�GCL�!�~~�c����L�)̤!�B����!� �j(d����?��-|]���1���7���+ϚnlM(��̉CmC�;:w�e/��~Mׁ0�ۮ�/unq�\����a9��6)Oh;r�H^��/��dρ�&��c��q	G�/�
-o�A��(b�'�����p�"�N1�J��nԠ]����!y��&,�z�R�Hl�&���V�<1Lx%y����Pk��ZrL��wb�oz��c8�ϊ	�>ޗ�!mF���Ml��`7���'B8����lvf݈�{��Iq/`l[k�cNH{f��u��_�'�8 �;�Ly��D{�\���9Ґ�e塭5ڞF�<2A.����7�Ԡ��3-i$��[¿�	��YV�/���@������A������ui��ّ;��g��D�Mƍ����\�����c�Ϲ��߶�P�?y��˴�.�1S��<��F���5���W�^mV̚Odw����2-Q��p�Ih^Bd^�$���$�~�"�Y)5ѓ:t�h1�*��H�p�mQ�n�}@�v&�Չ�jtd>&�,!3�z�apH@P�F$i'6�e�@�GogH����I�;�`qz��y=]2b��fa݁��~�$����n��P`V����J:j��Ǵ�nbP��|�����L�@C}�e�DV��קf�k�!"�y2�՛K�u��0^/a0T%y�7��:@fu^w�
�.�Y�������Nu)�>B�;l�V��t<�B�K�3!��/II� �].�8�.�FA���N+��&�#�\I�~�"���H9G��h���#�/�qu�fu�ܨ�#/�kz8:U���)�L"��"�-��=M14G��e�p���CU���Uu~�H�-�Ԭ���r�	GEM#���#8G}� �k�����'/�|1s���h��r��*�$��	��(���%|q3�9V�{�x��{"��ɔ6�}����<4��T�F��B�hK�������ȏ�Ν���Auܷ����j��ޓm!�$=���^�'{�3�-��;q���G�p��W������npϢ���Vn�m+�B���hiS$ϛT�v(���R��!M}iT��*�8�-��IC���X�[��W��J�f`�9����ʊ�BҍfQ#�0�K��2[KK�4�)m�੯'�s��3�ι�����1n���ҩ�sK�,��X�}n�؍|��x�<�.�g�"ZD�p��А�Վ�ېJȧ������h���c��e� ��{ ��*A�9��/?�����`-.W�
#�}
s\�m������1�36�(��	��=����w�3�L��)����<?��d�bʙtY
��!�UC:����f�L�̙��0J�U<��V$㝈Ŭ�;���%H��@�;#B=+����+U�&��%�{Z��n`d,�R/��g��	b�=hҽ��ݰ��тS�������(�I�R=�6_�MJ61����Ȱvp�z�l@l;~ �WX�Y�'����`���տ}�puu��a��<���ei)�G��P��,������!��G�PDd)��[�r\b�>j�)�H(]9���.��֚�_J>og���]�*=����s�vl�+t�[E����ܛT���K��4@���I�PJ��|�g��#��Bm�����b����+��zޭ%k�WY{@4���1t�Ԡ����Xxh��|CC騄���!��<A6/u�ȑVAѳ]���b��sRj!�C��Y��nɀ�`�hY�Li����Y�$p�<��5B�_HO� Z���?����u����ai���Ą��� �EzRgv	�5k����|0�E��������t�8�0v�!6T{�uv�x���~T_(��v����`�VB�|�3��j�aO���� �]0 %_!*0-��D��c7$���
�B��, <߂ceRb�3Tv,�J�����.ZE0-����"��1����#��W!��]���~���<�R��*�LA�i�_��-=.Eۂ:��R����h}�}td;����d�I��>��	������[��Y�g�b��k1)m*���i�<ǭ�'*0��b���Tz��&��Y"m�k�d��uMl?N�J?�b�����{�r��Ԯ�\��������Vm+S��[V:h/���Hl�C�Dt�
+��K��Il����N �6��$��h
x��=1�*d��/鲣�P=#�%���4ߴ'��%2����V�Ỏ�ДY"���>�����"��v���LJ�\;	2�!_�j���+��s���9�Im�L?l�Z��I7o��?~�U4z�.SCz�r�\<kzd���#�A�,�F��9���JMM�����t����o3w��X#i���Ga[�?zZ�V̾�n{��s��DD1��K��@ ��<q~�������V_�v��^㤰���fy��k����u�������'֕$���c�ͷ���g�
\��ܟ����^BL�$�.ax2{)^��#7'��-hr�ߵk�J��|�z�!b=�ʊ������D�A�`�z -��Y��\$k�ų�~��Lw�$�"f:�4�U/ͿO��JDW�e���'L{��$$�,==i��jǩ~� �a�2F�m�_����=-�y��|��Ӌ��o�G
U����P�C@จ��o<����U��[y�U|,N`D&k�Q�е�̢�&��̓ˡ�����{ɭkZ� ��w��%���P�S�l��h�����\|�����1J`��C�o���޽��^]�����LAC�&$�+�7�����;��԰�As"���=3�"��U�"�/"�"3E�"S���B�A���Z4��KT"cPź�_#�Z�Y���C�p�L�wӽ#S@K�Τ��N��� W�P[7���!�������Z��C_텍�g�J �*�Ny"wЊ~��>&p�b��M��[y��Y���S�Y=o�zk?�3��������j)��ﳤ{�T�v<|��Hs#�A��#=��cd�Kn{���wĢ����aYkc����*)3;az��3��N�&��V���3�g�(���R�DY�<�j�J��ˤ���̍�F�ƭ0,S���X���A[����Y�m�v����ۧꨓbm2mW^s~��0�ۄ���`C��|���9�}��'�})�|`�P�!)��v��,8[�s�W���\�QF9�P��Bx
�!�^�.�XI�K�����q���I`�����_@5�L/R�ۭP�4���--���CJyE��>Q����#G']�:ZEc}���8���1�;�p�6�'r�JP ��$��:4�y�r�1���fLS}}`/E1�A���AA^?:: �y���^��a`����ɞ2�w����h�؀78յs�����팘^��2n�^��$i{��^A�������A�qY�]���6L"|��K���G�OS���lے��#5XNl5��޽{�b�x��&�Ǝ���w���]�X�_��R�D��$=��g���"��$r�[Q���z�K�jMK��	e��q�Y2�9o�<{O<��"�=K1�H�����E�e"?���[����٤�S%
�d:�S1�Od^�x�a(��U�ۖNOYEf��!jc����Rm�"d�1�o*�@^�uH�~��i�<�j���7�m������39f��Q7B���9�<F�5ՙ?S��2N�O�b�5onwf�C�,QoݫH�!�0�l��i�ɣ�}ן�z����lTd� �?ծ��D�������υҷ|S���}Ə !}�p��D���vi@oS�~��)� (c�~T"b�?�	�7mڴb���bF��e=P�bW~�e�zm�����Bz��(l�@��l,���H��l608S`�V�����4�D�7�0����C�d����K�����C;)��%;�����ߥ����\.���*��u&�J$�԰��'����_0��sK�~;Cq��f�?Կ�������23Ť�ِ���]�ic����󕞹@d�%�RO$���3������=-��'�b����j˨�(������"|^����|���-���y�砯<+�:&�j�*��������������3^M�'�If!ũ�~�!=��KC�$��xUm�VL���!A������b0i´؃���[B(%� ~�Xob#�Q�u��̩���,"fB�se��4������&�
c�^���=딏����W'�_�d�P�7�evD��N��<����EGH��Ԏ�~O��i�rAt��'�&��x`~c�{t7~��z�3��~�|T�.k?D��7��n�r����g�crp�!H����-�I-�[ๆ_����7��z? �\t��xlHu�h65!K��<E�_yz�#�^�ٴ����"�P'�h��,-U�>��a�~A`βr�txl�	�~�4@����F/���$��]�Ł�ԡqb�������({"� ?<g4�S|���¼A偅�����qu7�N���S�:�Ȝ���)�х�~�X巷���sfe�^�c���?���l�����˭D7l/�쎚�d�_.��ߩ�s}sV0���tj�P�)jz-��������~ ��.��A�]�R]z�\g��+] ���p�<��|
B��]��.��s����SdG���'U��r~���"ks�%����A/Ÿ����<H��]��4}��:������
��5��8CZ���3p�r�?���tK~f���EO�o���Ȫ��-��}�%���ƻ��ԺsC<����Θ��'����I+o��1�qo�2��"�.�ųH�[<��	,�8N��K����!ĉ�֏����v�8��(�����#Ky`d�����u�*ю�������s�q�� XI����p=�&f1�cG�(��*�5�e�����r�ܒy@oUѦ�#�Q�>����BQM�����FԶ,˺3��N_�O/ ֔���ݑY,-)\�hJ��rj��=,�'�ߎ�$`Y���o�_�>߬D�:��*$a+�?�E����$_.�1�v-`0�V�����Tk���xv|H�`N�n�\�^̑�s����%��w!tB]5�������f��l@�b~'����ru��ˆ�v���2���C����3Z���ѥ�u��>��է�r '����-�b�)]&��`��:�xS�.l8�y�T��w#��1����g����ͅ)gMA3Q�a�fQ�{�P����zg��6���� ��l� ����h1�N8pqp�����a�杻v=�c�.���a#��w˻�SR���ּNM� 6�d��"�}ҟ[;�-�V%<�<?HsL�5�0�?tǺӝw \(������G�r	#���ϟFcŨZ���e�-U=C�H��Nk��.�e�7u�̳C+�����u��������5�=���L�Ѻ�X���#G��	A�۠�xBU]����1�>M��<�Q(z��$"ڱ1|X8Zo���]��ps�MT����9z\�v-d9�А�N1h�R�	�P����<J���q�=�
�N����b{�%��!ێHKg��+��͛���f%������i|
R7{�����aZ���Di>W]�9�:��M��P�����Ԅ�ށ杮KF�]f�7�B��5�,��'ϋ��ģ\Jއt�L:��y�f�\�nQnn��2b�|����B��J4�c��p??�V��o/���hJ<�ߨ��wl d�nD3zb��x�֭[Co,�4���K44?Ɂ��0�D�{������S�\�ʯ��QA\�YHrU�[OX����~"�p��f���3��v_UoMT���� ��l���f55�Z��(��l�cJ��g�）�H����Kb ��*�}�������-|]�KI�&k�^�P(��*�������mC�SW(U���k� ���7�0���/@�KDv?u_ ��@�PtM��f��a�Y.Z�(��k/P�����Ϡ��p�9��I�9bJ��|�Z���l��	��4���scM�RH%��$�)0X�0�㲗=�gG�BG顤U�ӝ��h��N�%F�B�)��j�n���;f������`�ɬ�j:�;ml�w��򩻵��
󚆫+**4�lb�����T c�a#�A}7�r�0�͖�C.�Yw�ޭI,N�w����o���^|���?�V��HuA�iUY�'�6iū$���(��Y��Ь[]�:�ԋ�0�5�k�P����C�	�_��T	ވ��S��o�����Ϗ��8���2����tde���@WU��1-�cs�D��}��z�Λߡ�)9�%�71Z����"!�Y"��d/�V��]Ҕs��!w�<��_�1n�����e �\!m��QȨ��[!��	�	�Ro�>|�1�V�r|���ǌ�5����Ϛ�dee�!nQ8�Qq��0&S�-��e��D��n�52����l)��/��b��2V�l��P�M�C�����9[?/��X,^�Ou�c�{ޔވm<�޶��C�p%v��Jݞ�E�n����xb�VH���'o��tp��@���ng�|���.���n�أ�7��x ��x�-�����k���UN:Q����� ��7���R[I�1@Ԗ=��e�!�Re\�]
|s�ʃz��j��ё��ųS��4�R3�:�[-�(t�Z$v �����k�.Z�J���%��.��j���W�L2��Ԥ97n�:@�$�����Z�f��`qQ>����
�a<�iI��.�����~T�(y��� ��*��߹<����㍘��/�Txм掠�� "�)ڤ�x8���1B5�Zw���ˠ��Q���r����h�S�'v�$Y��W��\PP0��;x����2��E5����A}|����@�� ������u�qn��\<�)�a?Gy��c �t]��Q�D�l�e�-�~��rW�NޡE+�Ju���`�;����!�Y5��t;ā)XUB��Gr���%pÉ�#� �X�YoHߡ��S<��')�e4Y諌�������CS��duc,mx�;j�9r�#)�%���B��eD~u6]<�ooB[yV?A[�(s����� ��o�!�;v@8����`yRrl�;e�E�Z�8�f���P�C"}h�#;D��s?Fk,Y����w+66v�*��a��@CC�	�Ԡ/1-���UU�%�F\8�*�hS+��i�K�����������69ʫ�
<��A ߉2���6m�8��=���9�bJ3��&��xъ��@���Esk^"��Q9g3X�{rݖ0�ȘU�u�I�V̘6�(W�6�S��?-�٤ &����e�#2�#;��u��.ʮ U끠�)7c��/����}����������4����Ё�b���a�a'�vݘ��g���aa�(���tv�8�(�BT����0��D�w&������mp�����}ׄ�����P狁n��6V�ǜ�#�m�h��1���C���:㍑����x"����H�5�ږTP�9�ʸiݙ����#h <R)cz5a�����{b��.Yz�oò����z:F�LJ��7�Y�q'1�5h/�)rI�%����ץE�B��hMݩ��i<��6w��Yu$?m�����T���ߤF�3]d�D'��{���>��EM�P>Z��q!T�_�ñ�̊�<QT�*S�1�@���F��w� �o��2e�y���:
f6��ai5C���՞)X����H%H��|��3�mb|,ެ$	�\��4�A<���2�ʠ��Ϟ=���VhİO�=��w@L��?�+�m��D��,������H"��ug�I�5�J�v����CG�U�P���V��u��(k㯮!�Ɖ~�r�?!�Ӥ�m�b�����]�?ae��2�)��C��|��`b��xOHּp��N]�z�Çjݒ��3�@+�n�p���;;ZP�Wz��z�ׂ�O�d��\��(u?�˛)u�����첔�
X�������}f�
��v�.D�2B�_8CE"Qfy�'�Њ�ֶ�=򠪫�j!k�ۍ=�q{�(�*]%�(6ԡ=���{�c}���L�$�����&��ai��Ό���(�e}��zȝ��A��D}la
B�A��[A�%]FK��aЛ�i|�?�U�W�u�þc����A��:uDx'�cj�+�A�tY$�V��CFffx0XjՖr\�7�"䷌��%S��3#�#P�#�m����mN2�Tϸ�f(����g�m���L�1/SU+z{)*�7;]q]]�6hmI%���vG*T/���ˡ�K���H�+)#mV�5=m��Ѩ�H��nUi�l��ٌ���P�:֚y���IrCÄ�v�Z�SMAC2��Ua'�K2LJ, �ǉ�_CI�ɯ�z��:��:TmQ���J��BE�ж���iGQs��mݛ�Q��դm���(k�#��{��ŭ������j-�c�T뷸�U�_dRRK�{3�u�/�鮯)���6��ߒ�sH�[�x�ྜྷ��맮Xg�@����o��g+!�y���uG-
�>�!�1�K�%j��e�"�k o�'Q3��{��y��G�?"�����oZ�v�
��Ɛ�� ��JMK��^�7o^�9PzV�[���?\9,�����*����L?���פa��gcT(��g�V�׼�C�����.Doo��u��ug,]G�z�0��Z#��Ep��'��3aX���`���i�P!:�BF���:��(��jpʺs���̀��F1UH,�ynn�~֕	ԁ��Pw��*h�Y��16�H$�2z��R��c��S]N>���CI���^�q�����^�nC4G�lw-���1}���t�=���s�"�,9C���� ��5��<]6�UFk��,=iz�3�.���5ϵ+��
�U�6H)B���,�0�� ��EwI�Y�toB�9!}P�D�Q���U�އ�q܁)}E���RKgM���v`�؁s(B�}��W�E��*x����*�V�� ��1c��D��Cew^�;v��c$+ӓp]��E�x�4$��H���t+E���UZ�����"��ٿ%�w��N>Za��5 �H!����tz�II)pQ��΂�������U�?|-��Vs�0�Г�k_�X׆ҥ��:P��eR�y�h��Ћ�\�������Oz�|���?O��YJO�*�e����C+��r���<y�{EdO��a߲]�w����9)ݪ�� Wa�� ڒ�����3h��(���w��{�m���E۷2�ēP�v|�%�9����#Z}p�B(������7��f6m�QәF��R���N��N]�쨾lV�	~�r�r���T�0�������@t>��hŇ)7fݾ=<b
B��;i/݋��6�1�ڕ���߇Xw�-@c0���aF�x�V�����NO.굄RJͼf������Jn�����q����W�?^���jn}�GfHp�������@��wіn̬`�}���C������s��U��S�;�l��JW�j�i;�m�w/��55�Ӳ�2OpF�kb+g���4�6�-�V[�G��3�q���ÉG�Y��Y7��8�[�cI�>��H�v5��ܜ��
�<n��fp�ԝ�98�8ȝ݀O���d�O<>}�I�~�]���|�II(�k��6/7�?9�����MvM���@��}~���p�O���q�Ol7�%� �^;��S@CT^�:Q�
��7�\O�޷a4	�]GP~σ�ל.kP��W�~������Kb�"���6::ڳ<�=i��P���[D��j̄@��L��i�$7�Κx����V�,J;U�Z�(��!PVD	�w7M܂��xt
�ߘ�4X�6"�S_�})�b��5��J��J �*���b�R����)����T��ž�|�W�u��R��Z8k��H��WU���&MT���C+,����n��j�G/l4_�5��J�����2�	Ɣ�ָ��t�7��G �����ne려Zĸ~���!�L�F����������e&%��Etls5-(蕁��L�mڦM�R��',E��5�0Z��ɩ�?�=�u��2n �j���A]��E!��G�]~Yv~�������~wwwC�Gmj�T(�`���dH�b-
��ֈ��)�EB��}n�y�[��Z�h/�;��͘Z�6�;��:�+z
��RfۮP�P�_�^,c�A�
x��*�����xA�k,) ��E���>�m��e��S�Om�82V�����������F���0��{�w� -'l��ԉŅ��?�.%-�T�{�{S���GވBԍ��Z<��LJ�*�>vuJr)�x�/���ݻ`V���(I������|
��6wdk$I�zVƛ㬯"'gPvo	�N>��:�xiii�A�>A��:QX��X�h���d�4`Q���EY<&ވ#�})��0�L��؉�_�Q5�o3�IwI�h��͘�(à{P�z�uT2�Y/^С�I/�c�;�w�^��G��T_(K�%��{c��?�0��_W�^(~��A�����%�q*G��E�ˁ/���52af�C��9�����e؟"|�Ỿ�YؑJ#|,8W������'��ms-x�8$��r귁h�/Y����P����S��F �y$��OEn/�VV[����#��IC`����d&ɇf@9��H�~��h�öQۮ���΁R5�]b�3%��ۦ�c�ju^��Tߣ����]s}r��V|�䖋�:R��1�ut�9Ʀ���(uG<܋�m��th��:^@�:��b����~S���U>�܂c�s��Ռ0&n#��*�-�15(q������� Ӓ^<��U�I�)z�/�9�x�}rCSS�zEg�+CBD�ƩM�]�z5�ڵ`���u�
�o��Yˀ�j'�"�=ɳh�_{Y�G&�Ώg�v�♧]5v?i����q����[�Qs�{��ʶ��E������;ߧr����"�Î{�ά������_fݢ3���_�j�����]�q`��}Ng��+�/�R��<���ƒ{_��h5��j���8}.d5�(P�u����r��8冎k��na�0���s@��`;F%�ŅI[�4�eH/�����s�D�75@C�\$�3Z��T�<r��0,��Ra�fq�}�X,�d�:��6�U��|Ap�1� ڠi���!M�x�0�o��#�¨�.��}����5h��:F�-�{13��d�/$��By%�/�P�rL���E��;�,; ,B_��s��2�.0�	��a�	M�q��Dq�z(D�=a�Q�60)���&��]�Z����=���]��Dw���}\#��������+�j}C�?ѳX����C����������u/�{��:t@hܜ��;0��Q�^���*��W=��贺1>J�9�Ժ��0�Q<Hd���3�OŻ}�U!99�<����('JU���{|||���e!���a����J�)/x:mI��I�z\���9ja�� O�P����gόc-��2�QV���o�)�]?�݉�V=���M�5 1u���L	#�Ip�$�� �8� k��O7����ar���@��OBnS�#��8W5-�ka���a��X��T\�,���l�blw3�0���)��:|��,����]�z}S(��ߢ�5Ƽq�[�9������(�e}����)�g������}QSq���{n9��ȸ��(�@ʯ���"��|�C�71�V	�`���7�?�m�\^��S$��5|b-�Fޜ�z��3�������| ����WGa��d�7v��"�,ժ����Ng�fv@�x��%�6݌����
v��e�C!~Ѡ�	e�# �Bk�9'��D��vI�����
*rp����`d��7Gu�P�d���=euHS\���N:�b��g�61�LJ��X�"�"d�)!YK�>.���Q8۬]̶Ԯ�T7����K�+��)��0�C(��r����EЧ���6S+0B�N�Ѧ��K� k2dl���������*���'��a�Wa�/W�}���R]���u`�/F� )��O�r^8����gڢ����f5��e(@B'�x	v(�Λڟ����ݵ6�*V_�?8x���T0���yi�����o��
��y���y��+;��G/�v�:�L��k�Ǣ��������{ø�8��\�����@�����k`������'������*�Er�w���՗K	 S����sZ��E�rsv�6B��!�"��C+55�(�|�L�(���o���-��w��r%^��2�F��_��4�K��@+�c8r���|z�]_-ڴH����Xͳ8�_�o"�����Q��20�7��g��w��2�F�SN��0������nb�T��'Х����a�y�j��V�u['�r%�\n��P>��d�� '����#L��Cv��4ۣP��Po퀝�����u8��-���Ŀ0'��47��y�r(��6�z׮�-�R��j�dqMP�L��t���*�=˞�(��t����1f%���샵�Vk �S�h��eee/C�����VP�Xa
0D��8����vΐ��c�o��S��u�j��r�@�?>�T��O����#����7X���ao9螺?�V�J�DO�c(�7��W�S�̀�ĉ٦N�F��ns]����6��d�Yǂa��������%��'����+���R�D����$G$�WX=��wW���)P'!��N�/�}؀J�����E ƒ).�ʆLo�&�.�
���}�ԗŹ�/�7�=�OL/W���R�5'�������.�u)U�� �zv��17�/���ۦSǓh�?Kr3!�籟��~���wa��"�d�Z��6�7��}�;�1*������|3[���ޖ��S�'�LA�����9Cl������T���v�L�)n���#��v��O�:]f
���6�E�}�>lt�b���y^%B̒����\�e#��c�Ae��������\]T�H�_�����[��ݻs֮I��ܦQyMŻѯ�p�r��}�	GJO�1j�窤��
��"�����������+���̢��6aڌ�+�J��>�h�H��ԗWoڴis��3��~>P��0C(.�O��F܍Rbr����%ɚ>��غ��!�[kS�8��%-��u,V����X�.����8�)8�ywC�e�e�� �GP.��;T_ҵ��-�K���6�O�M��S��c�p ��|��q]��� D���}��9�]R~!�e]�͚������m�q��&[�?:��� PK   G�rZ�mg��S �S /   images/84f81591-1534-4849-82f2-ec60ac1f84b4.png c@���PNG

   IHDR  �     �a   gAMA  ���a   	pHYs  t  t�fx  ��IDATx��ٮdKv�b��sNխ{ow��C�8u�-�����,� Àa���f�_�1�'ï~� �	�Q�I�I�d��d����V�9��w8��"v�!3�9u�:׽Y's+�5Ǌ� ��.p��a�����%'�x��3�z���K_/���SS�
�&��4-l6��������i\x���Á�m+��~w]>=\d�\�Ho���ү��k�n�t������N�5�s��1��>>q�>��ϡ؇�����i�&|B]��k�_�f��Ox����~�Wa3�z�/����X
8��N�C� <I�i�wf\=16�\����C�!�ZbN�=	�(L	�H�����S�q!����L��ǏV�։0����D��C=��VjS�@Ҳ\��>�޽��y�"�8�08QX�J��.p�<0R�������2/綢����?L�\d��?�ׂ\� �r��5��m�ٞ�.p��q�Ĕ�U�ѦK��`f���S�Bj��c	�~����U�;1-6�v�89��K">2���.p�\�~�]M��Bz��k�gk����Q�f�,�Sް*K��>��2�V�5<��&����jt$���R�B�����V|/����u@� ��l6-�9m�-��] �.4n�n��:�	���Ǔ���'ID�, S�2/�`�����u�\���0�&�
�t�琩4��WT�.z5�Ӳ���#�ѣ���OO�X���6��n���Ol<kk��q�ȼ| ���@@������	<�y��.l7W����ի��2|���p�B��V��ɻpБQi2'�%3�kʸ�N�t��.p�<��4/�������*�{�@4��gyG&?@���^(�?{�.|����\x��a��W/_���5��\�o�b�"4��9W�Y�G�k��f����;x�=�/��%������O�������;p���|����?�?���;߂��U`f{蚞z9�rd�ɫ�F��E��-_���}W��]���p�1z��4.@%��M��c,	\�XJ�e�M5�y�'���4�Z���ڦ%Ɩ
����ٷu8������<���������~�Y����ᓏ>�o�����=��!��Z8�;%0/Q hĢ7����О�"�;��W~�k�_������O��B׆�P��6p�����>����o�����+|��B�}w�vAs��CԾ|$�Z_��E��6H��L�5���E�%�rט��Kɖk�\�8R@��# �b�o���g~O�§��׶�����i��c����ƿ���|����=����߅�&0�'�`��K������v�������|��~�1�MÌtT=��R���ҡ��wۧ��_�U����_��"���P8c`�����>pG?پ?������?�����ß���p{��-���%�~�7�I�0O��S#�:�^�j9
j*����o�8��i�����0�\���x0���)\~�ْ��T���h��7�K���_��o��F梂<�D���m`^?������������W��W}
�U��-ս�������_�5��{���O�	����>��k$@������LĶo������~f�.<yzŎ���y��t̄��+�h�<���?�����������d����Kjc`oR$�s�	�����:	�?��<Zbl��K��'�c�����΃�]�0x��uS�F)�R����(�� ���H�	N�h�����������~����H7�w�u���r���l��Y��{?����	��[�	��p�������E�xb�g>�9���~�'��B�h$��t��i��~��g �N�ʗ	���>�O^}�6Kه�Hͯu3H��c�tPy3rK6b��A�w�;��d��K�<�)��A����	��!�� �k�]jI��m>b�4
d��>��t( �*Φ�`���B����_������I�!�A-Mb��f�fz4����ޯ�m��o���9#�f��CU�'�������>���A���PF%>}�	��W���7����V�+6�e��_Hᗏ�?�]c���A��4��	˼.p�\`jL�����@!5/
qߴm��@�זZ��9��z��W��/}>��/ �hM�ʊF]���Z��_�
l~��m�>��&DT7��w��wߣ�F��i��@�����ޅ���l`z��5�M�m���Co޶�jd1�����
�TP�0�sa�)v��^L�1�����&I&�]��� H��
��j��j�
�an����C2���|��Ablha��;��;����M��>C�q��As����Ce|�Gb�	���kx��)��Wh��|X8r���eLV��6I�I�L�S#��0]���A ��E	&�y52)h?]O!�(`_��PB�#��u�\�$����%�x�a��1����=�4�{�G��>�^I��W�9/��'�RBg4+fkl�ׁܴFn8�#pp<?kZ'u6ۖ|^X���?����Ls7�D̦,/�I�z4��m��nV/�����QI��S�&�C�:}P�kg^�8�@�2Z���pP�;��-���(��q���.p�\`!���t���ԍ�01I�K���Om$\��0skQǴQ����_'Xty��F��i�BӒ!/���'��pR'�,����>�t)Uͧt�"LT7���<��S��_}v�~�l�9�P	����9���1,��<�	�=/��\�i�c��F����$�eσ���߇�qc�f�H��vy�\�-�_�YI�򨩏�	��@�h���y	�dr�㡕�y���*�M/rR�[��KJ�̛��䄶��1{n��I��G�(���b�E�#��?�o}�[p��oZ�a��������t7?��7�	�?}.6Så���_����(�l����`4�#v��E�4$��A�as@��R�w	���.p/���X������yvg0sj0�m�40�m�rv`|]]�" o�9bw���} ?���g�_��hp+j ����N��?�Ɵ�?���=q,J(,V��jJ��اϟ�w~�=�h�)<{��d#&�'?��Xd�5�6��:�����G�����}�j�`�Ԏh�\8"'C%F&��2=�$y,��u��z���']�" Q���Ͼ���~�\�s��>��GK%�E/���rf%��F�r�$�U����!�L��1"�B�g"�����������˟� �R��F��؆��>�!�_������+�8J+eۼɣ�1��{��o�9��?�g����WA|ym���\?�».p�]@���k�i~�ۿ���?�Kxu�2���xox�@y�BƗib���갩T�o:���X)`C�LA�?i8�s��=]��=um��R0H��@+s��P_յ���<��lV�!��O9�|���NmXim�Y��Kxk�IA�{/tK�|=�"�ҰDa鳌�mtGEZ�K�5��`T�����my��.�T�������>���s?���	�����]`��=v��p�=���/����)�GL��{h	Ã.}����1�P؋����{�<����ʯ�O}�����h7����*�u���/>��O��7�����a���Γ��z������>�m�(Ih�@5o2m�d�>m�>�Joj�F=�s��k��[Z��]φ5����+�x,x,�IԆR=�l�Cf�	�أ�}bh�P�(��j}��U�G��4���WA����G�	L�7~�o�׾��p�dKL�ŋ��\]�6�k���{���?���6N4/���HKC+`+�6�v/����������?��������_��~�৾���\�ݫ[����Ͼ�u�7�'����%�����b���*���{���.ׄ�������Q2r>>�c���r��.p�� 
׉ i��՞H�:�w���4v��Z�f��%�J�k�{vf�3|2	er�x���#��?����߇?���W������S0��%|����[�]��?�7�G��:|J1�|d��mЕ�LLNm΂8z٧��=Fх'>~�)|�����P�������'O(��ڿ|�>��c���?��o7O�R�^�Y.���[C�+���7�ߚ����B1H:	�y�5.P?����U8F�H^c�ǣydK�-g%��
PF9��Y���?��c��A��q�d.��p1�P��FB��`�Q�Q8F��R����3������Bu� �����>T�	/���|������ѳ�'Ĝ�C��>��~��G�q�#p�۸��2��G�ـ�az�(�������~�=�~Ȝ0#��ǡ� �[�K�y��雤z�1' ��������#��lA��[g< �NMⴁ���?�t?�����dr�64�MLL��;Z��5E�������c���f�ǆOsB9�j����|6>��SqY�N��k�����2���;?�;Z���h2�>�Ctu4�Pk�k����7<(b�jf����vs���<W��P|f6�yq[N�޻���-<
�^��|_p`7F �q<�����4�@ާP|����r�(�z��-�pL��qv>J�8�LZViw�Z܄�^o���I��!��C�V�C�&�r���'b���lxP�P4��釛�D��g�#L��1I�� ��8f�i�X�ǂ�q �d}꠴����x���фce|
�>Eٮ�O'�kU|,���Ʉ�Q�S��CUdk��˱s�⤿�>�ݍR���D��˖d�f$B7p��w}��J?H�y>W�	yB
y��d�T8�rő���#k�4堉��4g��+r���t| f��dH�P|'�($�=3��q�kc6�z
j�䳑�敚�pD�,9_f�0���-}VN�L�Q&�l���NM�'��%0�Fܷ�	B^8d?C��'��U�����t��Y�gq�|%�ee�)Ô��L��������C�SG������7>p��Z�G����Q���9[������OFX �<v�a��Ō��A-C}�ʧ��������5�@��zC׵�{N'�*Ѡ1�ǥ�����)�&���t&XL0��%���z�۱���V���[�.���7�Ș�,�0�eb��帎vH��Jy/�.���Li�t��2�ҡv�{3��=e)y	.N0�^HW��t���9�����f�"�ZY+�*v�]ҍ��%![%29b
#�p�勣^h��]xK�I�n5|ļ���/+n�7�N;Kb9��c��W��T|���?KpI8y��r�X|t.�x'����[�8|ŗ�)6圊���;u���9��b|D���YK����'| ��19����R�4{��>(�c��{��0�%(k@����^H5kj'e��i��iC���S�����k\��������8�l�߀(c�k4�����/�,9�0j��M�6A� ��1/���:r�.oukZ�c�r[��EI��|��Ù��/�~p�2��=��b�JZ�8�h����M���gmS�2������>�RY��`e�W��ݵ� ���k<�y6��/��O1��,|��*���lm�&�Q�c��տ^|���>�G��,)'����o�1E�7���~�^)��@������V){�a�鿲5)Q|B�3�G����'!t���=�IxuZiЅc-�7:�f ���ް���fg0����S��#yFS�8�O'�N����Q�Rɓ.t���}� s��<��C���|l�s�R���RY�,���x��n/m�A�V��n��ʻ�;2ҦW��h}��K���t`���l�.hQ6�}�e��ӛrj0VN�Kc�aI0���Ɗ�tp>Za��4I���].�&˱"R�g4>�eZN�w4��,s>�����`�c�1c&�t������}�����R�>�|��{*o>�ܱ��O1���'�-/k�/[�7ъOO�a�M�h(��'Ĭ�Wb���5:�$Э� �!����bbX��-��B�(JҲ��c?[�h�"�λ�e+0Т'�����3�V�`8z�"{��O��������5 ���B��9��\�x"��\�٦�~����!}�7��o��0t�-3�C`|�H
�����0 ������5'�d�+W��8 �-�BT��21؞�;��v�YI���4��б����g���>�\��'ZN��.��N�u�4��`���4�$1>9Z�V�g
�%���Y�|��G�����=�,'�E	}7�O�D+�,�'��z9(l�Q�o�hfZV�5#Y|��s>.��y׻��A*M��a7y5�e��*0��:x�h\xi��H��D��J^N8!>�	mfZ�� �F&eH�)��G+�P�ZW�ا��7Ϟ��ϼ��n8߼�Y�F$
K�O��O�-�������h
KJ��ĖW4�
�Q��4�����U�l^������2��$�W:	b`�"�G��Ou�!:s=�Ajq�x�3z�$7��>���b��6H2<hW�6<�۷��b���Ah`��rS����b`�"_#;��(ˉW���0>�1��ߵ���[uFX�g�Hs��S�����5���0��8��'���:SNFXt�L-XI�Lj<�����̗S��̝��hYck˓�í���x�c�I��t���z��n7|	2/8xJ�o�ۅL�=��c�^�Pt�m��{��"�#B&!92�f���ˑ?8"��q�w���Ӗ���Z��"Ԋ 
�1��C)�k<�L�O�⎉6I��'=Yj�'��r��m���;)�'"�Y,T
�����KLͶ;f`�r(�.�h#Ɲ�ێ�_]דJNXu{��?�*�c�>�!���Pc`�$5��|7|tط�o��w�ob�����)�8W���1y)>f�>>SѩU|���6z'�T���5��I�@����ekuP��*+��_��|���3�?���=wj������|�L՜;���a>��Y�J������G��r�7L��quFf������^��ydo]�\2��3�rl��pv�4t���"c��������-��!�Kq�p �r��{�����3,]�K��WB�D��D�.H�hq�7��u��>���U`� At�t$��e���XkW��J�H���o�ɣ�_����9�@��T"�\������[��;��ބa�v瘹�
�-�c7x
�c�X�Ќxn�^���,�Y\>1`|�yp�����O�W�霉��H�+#��c4��G�-��q�3��"�A�,����:�O��Zq*��ӑ[Ҹ�yu��N�  a[�tA�������hJo�ya��ZSrED�e���n&b`b�ؑ��1��g��o{
0ff��_�{���s��c0``��E>�_x�E�4hf�&l)��XކN����,��C�����'	ı�e+�m��}:�)�.p���s���x*h|��C`��m��z�^�x̌�w����l�����4���gY\������ߊwk�ћ �L����qS3�-��ȼ���g��#7��i|��-�'g<c7kC�츇b�D*GFN���=dR�`�62(������	L��p0=����^J|��0ݩr[�LV��g].�$W/ۢ<3�v>�Ai�
� �aV|g�`��K���aa+@ڞ��\,�ex��]`;G�B#��t�j0���s��r�).�0� ���-{�h0�)��l2SPtn���q�FؠIC�0�
G=��������a/�d�O���ז�)�b:�_��MϷX��h��Ok��ⳤ�[|��Պ������������k|��§�=r��A1���#S������j(H �#�^� w�̩�>|�;VjȆֵ^�5C0͛݇�a&V�c>��R�*[��T�n�>������PO`�#�7s>�00��ĈEad2�}���Χ�j�eH�M�0k���ꢳ�Ďp�V�����D�r�4ppn�?���³x$�~w'��P����f�i9;�]�(]ә�Y,���,2��6�O-Xq�M<�,z�Tv6>���=�32�&>�����׃�S���2�3�s�q7Q�b|=�𡹼>��(�l �L�Cޔ���~�݊����~��.�-lo���Ag�@�h���SF
��*����|H��T�8i���y)5,�)������\��`�.�M}\+��~@�D�'�R���L�꯺��2�z�d)+���A;MUlz���R|'�2��m`s�	\��u&�!0+�����W�fλ�11Ѯp_F�\]_QY>��/�r�� .�m6�[V����E�pT�,����!���2��*qa9��ұ������{�B|4�#���1�-�;�*R�6����q&�(�q�b|�X���6p�=%�m�jþ|�u9�]6<����i!W�R��CqM��ń�=d��;��1U�(s�F%[x�5�|�cv<���p��rSB�vDU�t��di����9�CFh�ze_�k�nQsR�v���UЖ�[��H;'��_h�ю&��j777��
�c��O���1��
כ�3��SJA}g>:ݟ=}�7:W���Ȁk��e�,�Jȥ�������R����|��2�ۻ�d���K6�iD?0AB�Y+6$<o$�OK~h��}^�|A�4�%W	GT󙋐� ��}.�����ЍŨ�܅��gO���`sS:�۫[��Q�}҉���yE�Ǎ�I_�'�c�O�nB�$�5�(�O�z@3u��i�Vv���u�q�'�	=�xl�k�;8	nn���]��/� SV�%j0;7��MP�{1��r�*1�u&���0��mt�����n����\��<̳�G�\z�%���,��p��wޡ�Ѻ��)"<}��,Jw���4ﱓ��uW�ʱ�('"��ɞ�&�ٝZ6�f)������^�#���*e�c%R�f�y�����p�rq$����$�]~De�7���=�C<�%SU�-�K��� �9�,|=lR]<6������HD��a�ia����~>5�&���l��h�,+�R�r����540M��&MU�
^�F��,�Q��Z s�d��7X��/%kPC�[�T�>�Cz�<R��锚�BwA�Đi"�D��f͖Lk�������ˌF�f�͟K'W�Ba"�00�s\E.�3�4ݦxLG�Ӌ�{x�# �^��0nn���%��@��Q��()�.L�zJ'E�������oL�~�Xu��|�\��uL�.&O��1'��ArF�)�1�<yJd��?��Q��h�����8���E:ě��ڒ]k�Ӗ-���2
��c��kY����-nh�L�,�2X7��������M�%�#���Y�Q)ꊬ����2�4()hz*}����\>w02-4)"C�%!�<XV׉z�n>�ށ�NRce�p���E���|8������=$%�����h2��/_ҳx�?�)���7��k�ۓu	i�^SWb`���ЬI��)z�e��ߣ���Q��c��\����S���џBjs
=�(�˞����X'L��z����9"�bB�N4��v�S�9	��E�G[4|�5ϡ�*�8�5�R��40��pʵ�('W��.p�7�[�.�ߓ �W5�XGAd�
�Mr��WWW1�C(2�@���aY�W�k�[&��#w�y϶�$�V6�1�B�%Z�ڶ�HϤ��8�������o\t��u"�0m�tR���%uXbjK޵�L�QÎD&��P�Ζ�2kt��7.��jE�����!�s�e;�]��\4!&u�IȾ�Ԍ�;���6�1idk��5����֘_𙆵�9V�gv�w��)�B�B���5]���e�R� %�yr#Q�t<�BP�N	ra;1;��50���-�����2��n)�;2/}�=�
�����C!^_��E����ʑ%���
	��tލ�����8 8I��C�R��9ۮ�&(�����N,��!ҥ�*��J<����i����L��k|��a|��Ŕ	[>������1��a��H����|�)3j7���QM2�z���<�������Ͷ�g�g&D=i4d�����3W
�Fy��eY]_a�b�rm���K+��*^+f��ϾImV��Od?��z[S�tޡ;Ї��F
B[�7�|](���t
�@��50�|Rew�4���&��`�����֐Z�j��iXe������N� ��U��j\#�m�r.�$d2��@M��:I�XoZb4)wkC�V�v��#�a�ͻjB� ��S�9���#��\�TSvπ��.�Y��6w-՝��޼2���^X	}ũ"m{�/��b&��èK� N�FϜF���4et@r��	�I����Lc6,��|�Z���1�"�z[!�i-�B���V��?�������W����!LV��k�֚Ь=�rK�� `�^K�����%S�hh���Q��y��T(
���ܣi��Ŧx%Ze�:Y�$uϵø�#rC&U´�Pءl����k�2���(��,G�G�4E� \�Q�Ht�4ꆜ�-��h�S�	�O��,/O$\|R�th����!Zk������Q�D�<�x�ծ�Z��rV��Ǉ�_e�����_Gc>� c
L	��M:̖43=�9�n�A<AC-}���,� lT���?�S�wQ; to�$L�]0/ˬ|�����P�ܖcm�|�B���x��q���\��œ�'E�i(.(����76KeR淯�oMM��V��� ���|P&gL�ׂrV���7�Ϛ}���`c��ѵ|>�BY�G����0�,����dY��{6-���{`�^�
S)�{���"�������M�X)����g<f�������->I�$؂���&��Kҙ˵�R��|0�����S`��!FH�=b�{�̔4Q��1E-x�l������z���7�)���V�xo%>��si"]��jBm��1��������bT�5�;#^Q��s$kXO���<6���_���kQ1
.$��o+10%���7���X0o*�Ja�9��M�D�x0�ڙy���w�O����K�ٻ��7���¬�����?��������`-��,>��Y�ɻ~	J=���<1Y���=��ۂv?6|��R�Q��5Ж��P�nʁ�����j�K�~*/{S�Wq����&_3�"�<���\H�,��U��1b���0�]ރ�w^'�����#?�+j`��h ��f��q0s��(���(�.eqfջ�]껸Y�G�j��S$�58Fi>?��������F��jn�ܠof(�=Xf*[@���axt�,�7��x�#+�l%|����:c�7����TM��Wd:��uQ����A���.i�����<ɺA�g�h<@��IV53e-WF�_ԁ%Ӳ�s����b���;�|�b?���g\bb.�<i�tc���ʶd��"m4�a�b�ti�6&��g���IX���
�
�,������li��d�KJz��YTQ�2�Ķ�扷�0��}^��	�݅��s��Zy\�Z�W�wH`����i�d$4Q�9�	E�U�Q;\,[�6x0F��2SQ�t���Ati�eC>�ɣr��E�5�$gT�b�B�-e�h`�vbgLN|��-M<\���y? ���ٜ���O�I|�kb�G�c-��>�u:����T�����}���T&Fځ̊2ō����n_Qd�v�$VS�陇*tgZN�Cfͅ�����z�w�ucj�ڴ]KX�X�1�Z����]���{c<1�R���7ʻ=���C)��q��ҿyp�{(�Dm�[Ɠ3g`��t��LҸ�Σ$�sgM̈́���#�\�h��o�e<���A�#J`��X�,�PJ�������-������d�B�)����ߢ�a�`� >�O���FR��^��2�T���r�Czާ��#^��4�}����-G��{���81��Gs L9V|^ڦ�����j;U�4t?�3X�CJ�ʏJ.��F��V���]K����QzH�{���q��,�`4�L��;XCy�``ŝ�މ]r�t<�t��q2>k�`���L�����_�8%\�m���K�����ᒄ�4�vM*E�|� V�U����:�>D>[֮6*<����$Б��Y��d�aRGsHO[�2�bR���b���䙙���`>c����	c�=��N��O+�>�ɴ�*�m���a������W��KCKmx����z��T���8DG�ln�1����eQn���ɔV�W�6<f|&�3��#����\<EJ�����Ȝ����|�k�M�yYg{���k�J�q��{:��5�ϩ�,M�-Z���PI��AVG8����A�>
HJ�Y W�gQA�U���$271TU�h���i�m���Ĕ=%A�^���{�1�u�an�UtC>.��}����`j����jI����2�7F�v��� �K^>>i@�D�����~G���m�KB�{ѶW�;*���.�X��x=$hu5�:�ъ]��Y��6��dy�̠��F�I��*o�FcH��c����ͅ��?�o&�PLj�>��\�Z��ր{a`.��N������r<6�-�@<��m�X�Gg�q�No��Yjf��&M���,�|��:k�TK�7W����h��3j��?=�?�|7:r�����f<K�}����p��=+Mn�T�h��_�w�&-�'kAS�3��u�q4Ϩ:�D��E��tJM�¼��<q���j󡸶��#��W����Km|0&�--(L��q**�u��2����M�ިi�=���m˄�ė}�1�%��[�T����2&)Wm�P,,k�[i���Hi��_xM�ǈ-�5G�@P�v�Dʙ�,8�ȺC�b��V�)
VE]�ۧ罽VH�z��Ԭ9�D�9������j�)���r�8�k�T	���c��^]�����|,\w��7�+9��J�D�������\��ά�5n���T�[2���t��x!�4哾x�+��~�00Μ��_L^�@<��8Mn�$cԸz/�N1-"��O�C𻆧vYx�18U��:h򍓠Ƭ�Y�N`��5�ր��X��O?�	8S�׺�0x�������ǝӾ�N7�{h6[���]jk�I��s�X�XNJ|M_dv�#,�\~�`p !}���b|��.C,���ն �ێK�o�b3 �
B ���,q�h��.$�<mƉn3��]��d����=@V�T��im�Ӧ/�1��Vn��l��٭��E|�
�?�~z=�MN=&T)б����P�\=�@;�6�����s���P"WT�ކ��i���A2Lw�i�=����Q�"}�BF =�Cf�-o:|J�TC�Y\L}U|I�B�ԫx��c�;�$3���#}����r.�V"1�3���r$)C`d(<!s�k���A	�F6�0���i�=��T����Uk�\�?��<����
>�ά�����S���Z�eo�E���I�X��5�e�dk+!��C,ޛͽ���Ǒ��v{�� ]ǩ�t�B�˧yۆy�J�D,R��o>��C/����W��O�V}Z��@f΁Rʲ,/�q���U1�$I�(����9#���C��s�:.MfFh$,�� *F�T*Z*F ��ʸh2��0�psaN���7�H��,8m	�C6�� e��I�D��f��2���t���O�T�P�-ق-q��>���@e��,bC�?i�a��,8�&#h�	������W�HfN��S��u������\�I��^�!�~Cϣ���!>�l�і�h���f�Ǩ�����ݛ�Jc�:�K+��(����q���W�GǛ�4DħY��0~ϔ,�4�('�1��r�?9>Ȕ��O������_��!�`�
Bo��5�I��#�cu����J��pu�^S��C�S���4���*�����v;����/���W�OC��7��-Mh��L�4����K;�o��l���0+]+��&a��yY|������8�yf-
Z�bV�䋚84�J<Y��ɀ�#0�J[al����N#���76WEY5G���Ag�؅gi`b����;_�T�D��4���1Y6�r�HOZ�@L�>ΔTf��g~�q!(�����C|8�)�˱�Ç�=?,�q[H� B7��$	o�����Ԏ~�����{�¼�������ߒ�uz�k�		2e`�Y��o��3�>��j�
lDϷ~̎�+���?m�\�ȼ �X%�t���П����7�s��2| "ð��O\�DF��̕�Sl����CBl�t�d��ѭ��=�RFK�to������a��iW�A���\�.�#@�7T���ڞ~�q����>N���'���l� ;��@[vD��O$��ܦ]2-�Ŧ�Ky���m�Gk`fsx)g�D�?َ)o�Ldb� Q���Y8e��N�F��̫���4!t.F/:�1��o�w:P�N}���n'�^�ER��μc��Ϫ������L̜O��&�{S]ݲ�dy:،gs���^�ⓗ3��.�P�M�=�O�x���&-�F�IĠ1�K�"���ِ�i`��,=����_����{
�O;٪�����U�p B�����?N�n����� ��'6���g5W:o�s2w�`�a�5�Ǜy���<Y�$>��6�DM|)>Y��ƴ�od%�1���i9�-���ޚ���U��):5h�8oZ������[��M�(�찿#�����w�n7c=�S}X��@3z���Q_�n�����$c��N�+�!D^$�%�̴��-�=/ú1�&g��ijh/ӹf.��%�U�,6�"S,�ɧx�ʸ|¡��w�ފ>0ь�=b"��5�ס�v�ɠ�@&,m�"�C]�t��d���0��yuW W���'��[;8
�]�:��8��y�!(��@�Hf�C%�D��r�ę`�����|
F�k����F��\|���Qg�2��Z��X20�,ʋ�䎳��ǅ�>����۠}5�k�k�uN?�&�d�����	һ�����b"9��+2�NMY�O��������#��ʵtϖ�c>�τ�a�ywp>��rJ|�)�-D�A^B�x�Xa��78u�s4�gp�cӓ5�[[�\bj^抣y&���&�Y��K�l/6�u����ۻ-�_Q8kה�Ǭ����M����*���Ey%B�� 'z����������d&�:�:���]�`Π�~�.��'1�I(���W����cmK51Ά J���2QB�7�g�oF�2�r04���u��ϷAҾ�7����૿�����s��p��������h^y��s"Oߜ�3��80?�/�I�X�t~'��Cl[N9}�#���/�������-�/F��97���!����0@��R�c�Q<�[�����$�&�U#ND_��������^̓�
C.]鋹��T2SS~&t	�p�O�42�$8�뮐�k!e� ��ׄ�,�o��0I����6��ږMꚂ�+�k4m30�F�2�
1P�ld���d0�����ǈ�e�g���gX���f�]��n�|��������o��_�f�14袑��"F������s�r��� �adW\[��xⲔ �&��'��ļx��HT�{ࣳ�@RRk����C��k��d�c�K�af��$F?�m`\���p�����}��l<G�Bɕ�M�ڍ�$�S�x9��r�X���O_{P|���x/�8����h\Z�Ȥ6��%x>0�z��	=���h��r�ɍ�L� C��>��fdȊ6��u������T|JY��/$n��t.$"��4���]�b_�1��<A��( ���%��5[�i�Q�Bc�{I���)�$�+�f�dZ5�Xw��kV�x��le��wp>��x��)�|�o�V�(�r,�jp�09��Ж`�-��\'FZ,��G�C�[.rz.=�D�����jcgm�	��02|E�`gJ5�jCA��PsA��z
$�:����o�D�ۥ}�Q8�&@�Y����B?g�� @�O0_�v*5�y|�͇�r�$P���g�q�?'�cߦ�]CF��
Ù�50���@'&��ֳ�ͣ�%7�A�ö]�A��ru���r�E�L�S)�`Rk�ݨ�QvE	���sY76G�l�9��M�RjU
S��ڐ�]i�^q^���PR�t��Z80��)�Eho�=�I��9q�b��&�!Љ��楝���Ŧگ��2�k�W�*��
���/ �ֵ����"s}>��P p泚�tP����g�F-==Ƃ�P��SIճ�%rC;6��;�Mӌ��m�8e��c���eWX�.��=����w�����'3!k{��!��f`�(N�_��!����:V�w���<�l���"�3���w��"8����P�9�����$��H��$��_��IA�}J'Qm��K���D b�����U!�1�W
)ؙk�xh����,�P�ļt6
t*����!�	�������Yh�f�!�<�
:�d��V�KQV*�&�tK�7�F4���mw��}l
~Cv�σ&����=�F%fL�ۊ�}h�-C��$�Aߖ�1�G$mLw������K@XmW�M��9;yP���|$7I���ר<
	����kd�Z=�T��hĎ�-g��m����X���N��^:ϪR���@L8�/��� �Mt��J9�,��M E:��^�B;�|LO������Es'{i�܉MV���E�&Թ:���i�m��)D7�x�@���X8��&�x+9#�;�!gB�c�t�v�!�q�pT��2O�ɦ��`����k��Ri�/��p�>FA2��8�-�p��J:��D����C��Ky#p<F���h)&K0e^��̖7�zv�w��E�bm
�#���*m;ˀ\�ʽ�x�åC0�j�C�Z�>G��~��(�����E�%�('ذ�� �0`-I/�:��|rfeT	ۦ�H���Y�K��8���4o���sj�x?�����ΕS���̢v+cyE�% �6J�Ԅ�%�����*S3�4F��v-��/�=S�m�N��ST3�+��MݪGy�����\��A},�t�������M�+�7����w1�Y�=��HS}��$���c����1$ ��1���G�-J��O+'/��{�\#�=�Lh��*�a�F�L���������h
�\��׉��/�d�&ל����;,mY�@�(S!'�����gNV�%����>e�q�U��~i��Vs��+��ꎚ}�g���N���M�<g2:�l��y��o�x��_�J�&��P6�ҤD�bˋ�d�`Xo&�9nS���Ř�ݖ��7$Gr���P�oa#ݼ!���M�Y��_���D�`�0-j',�E�2Ek�����D�(\��}�w�m���>	=�BF�6�a�����\ԭэ�X��*������K��g#��&�w@�N�G��?i����g�ѱD���2A���I]m�%��c��h^������>h`�&�0����륢2������|���$������XiX�] ͗��$�>M��rc�8�Q!��k��gT�4C-B����tp5�
[L�z�}'�5�|��)�U�\��b*�@�q�,����%�>"�/�[�As���I������F�D���� ��ƾж՞3Pg`�q޹MJZ�n:5�x#��`��,$�L���%Wb�/��Q�!t�&u��Ǆ	BN#�$σ���M�c�EK�$���1�O$yv*��_2W��g��/`@h��$h�(��儑�|�2��M�S�����T~W�hd^\����MV�į3T ��e+�259�Ks�ģ̶�r2�[@�G#ڸuH�W2�a^H4����YV0�Ŝa��S�\��}����p���C��!�Yj�rWT�O$VX�!	Ӱєv�1����(5o"��<�fx>���k{!
2�D����;(� �>VC}h���$��3�1~��c��a��_t7i+�|�ݞ������F�Wa̪ﲋ�ѥ�6�	�����-Ƿ$#3�̪ϳ.���q��|v����s(h��.�@5x�4g�;��<mM��W��>���$��n���Fc�E��4�C>9dIt�GR�Wuş�4G����91#�u��Z�-�e�Xp�b2�`G�M=<ۘ,�lk��Ad{dF��O��R�A�߀�z��&RH�3��<(;aXbV߅��?������~�K�Gӳoߖnø@��5H�����[nx���#�`��u�{�s��.	��t'D7Ȫ�m��tm���V��S��=Z�\�f[Pz�4�eť.JVJ2,Wm;Tڮ���{HqYE�EU��ol���=dHgm?���8;ji;�{(�ѥ�7M#SIr�l.���MYr�u}���1΍�19��Zl���0����nv1(��������F�w��^�XC��h���[eY��x�?2>T��_�=���[j���{�:�qY���f�G��<Rm�i_���P0���Q�_*�x�onS��:�
U-R*q���u�"Z��r����y4y�h�;�%eJ�ՙY�$�xMD5��{ ����[�H�G	fȎ{!�.j������$�{���������^���k7��+��ֱ#��'z��G]�)x=205R(����]b&�A����Fĳ{�����@��]n�s��C!搖�H���Ѫ鯅׽��h|��?�ͪg���9�y�,�(�yf�9�j8�I ������b���06�:"��[���x���,S���7��bs����><<��zk�f���L�(�}|�����I�	����������8�/�`�j��G�ػ��Z~��kn��9e��g��]鿂�f%�E�NKu˩�5�M=o���Ey[K��:F�ܜR��}|z'���	��7Ÿs���g.�:'��כ|3q�(4��b�s��}���W4�o���ńs�{!�Q�S�g���z��wA�5���V���sB��
������5�}��P��i&�fA�j$��T%Ӱo-(2��Ċ��f�:Hk`d^�Zj�k�Zd���ĉ�Ǡ�y�bшd�sz7o��$�_�`N� ֿ֕�B��F3ihx$oVƬ�N'�}:���f�e�P�,���(e&�$ ��i��+/1'��=^8�+�W~�����e�Hq��kn.��Pݖ���0`\K�9Fь����>�d^�z� �4�q�"0�g�������� M�_�lL���/n^�P?�
5�_
�����kI��29N��&��G�%-:#-ή�9-7Q�z��TW�8�r�ρ%xK�~�@���b��
C{��`he$�vC�B�{H{��wo����T35�S��o&h:'q������c�aM�=��ZT�̕���V3�����>�I�Q{��][�%�qrs�ߣ8���fg{ML�UI�~ +y��%���Q��L+�I��&�cE�ʕ�!��z��LO�9Q�۠��G_��D�M�?Ζ7�x��ϱ�	d-|�*Gh�pi2��ɵj;ԷO�9��Jo&������f�~���qS�q >�^42=h2s�x#�ZUE�]���U��s�b�]Y6�Ծ��|�e��2�?4`�H�"k�(Oj��!��2E|`%���I������WY:�l(����v5jO��3Ϧ�<�S��9_z`dor��| �=7�Ku��rܨ3�8|N.Ǭ^\i�:�֢"R|�� �`^��^�ӷ�y%(��M�f�����Y�8c+�'��%��)0>}�US��g�U7{�X(�2�:S���N�Z[���{n��t�U���`��x��0��Y�2�R��Q���k��Q�W�;�#���H.�cN7�s��F�G� ����}NY#�e���߷OL���`��YsOGɼ,w�5����ʪ[q�ٞW!�s�=�{4��Q!�ju��h��f��"$��E#^�ʠ�B��3������6����r�ы+Qe	�,:c���r�����Ɩcev�Gzs�&98��j�j�,�N70Tk���KJ����K!;��{x��a�ٴrd
�+>�舙��W> Y�?��OB�	pl.9�0#�=���N§��T9�!L+��e�E�|/��TdrOl��8R�1�����s���e�Mc��x}ꘐ��o��n����k����sm�n�Y���G��$0�囇�$*vn%�k<Q�<�n�s����z��ȋ���w>^�G�U�+ZXn��,-�����~y�\�	��~�[�
��"��z����9����^���/�kP)����a^���3���r,>産WXJ�����Fax�E"�R����vS���Hj>g4��d7���S!��+#03_Ts-^Z�G�7��!	V ���}m�~o��v�卶��^��皭46IO��E�e��MT�|�1T$5�w�4!�y��/���\A��L̛u���7F5� s���4--�tZ�Df)�u*c^S�	����p~�c�#eT���=��)O��]���_Z�x9����o��CO#K_}�����6sn�C�ǝ=����Ϋ��h£kW����d�~�;�QCκ�Rڂʔ��m$�0	3U�ճ�(�	�lN�]�^�c�\�' .J��w,�cRh܂1Ȣ�D���	�2=S{m�?R�D"�d��b�q�-�3 j�P�{��V�����[-kSbE�?���_b���C��7��M���(�=����nTvl�D�`�]E��P=�lx8��-�X3��J�w�8C�4*n����Ι�QoF�����C0�!����AZ?H}�1*�,�@t����T5G@2K�2��X�z��s=�c�U℩`n�F�߲17�̌�?��b�ۜ�yN�x��yu��Mύޭbwa`cPYкp�����5J$v#*$&f�Bt��EX�<�]hMC̩�>.�ُvq�P͇�B�M��v���Z%���lQ���&1]��1sl�gKHsUiq�\��)f�m7�݇a��\],O�l�%�4^��U6}�(\x��cm�Q1?*so��Ȉ+8f۹O俖�8��W�t.��@E;�N��F��;��<�ж1�����t��}\���^Z)k`�cuH��8;���]��U�;�}�._|����Z�f'���X�"��yȘU�[!�i���e�!�H�TV�lJ&���PMӆ�/����z>�;�/}�iaΩ �z����N�h�N�c�Y��"�H�©���L/��5#�ǘb�\�j����������1��T�78^׶�n��X��Z��"�'����e:S���KI^Y��/Ggi-�)�"�f�T[���F��yh�@�����E8̣DuB�_�0�JZ�U��˫�2_�]2,��-p��y��l�c~��Y�<���0��Je�):N'͔7�W
jaBO�A�u��j�1;�R����򕲏輒^uCin���u7�>�����б��Քi͇S�5�z-"p|>���f�]܎�m�*�0�I:��e4qa�f�9]�a*��XE���씅�7�^-
,�ȎRa��*�W���HS2Ov�2������w��j��a^�����Fe�����x)"�N�Q����Lb��	p�j�-��^�����Ke���cT��Z�[x�W)�����]�����J�������4~3�T�&��fT0��
��r*d��
ڝ0,6k��;O��(�v��eL�1v=%ƥd�jz�9q5B��qTSWN�IrM�s.���^����۰��~h%��
���{�<���@&Z������57�N���|�ZA�u]'J�?���#S}�T4�*����VU���L�uL$Q��7:�����f�^B�g��-^#���ZO�/�d�er�r�N�O�;8�,�%�3ѕ�������k��hW����E!�)x��Oύ�f��+�	��=��ʌ����K�E�>�����%10��Em��_<U��3~7�������?�vč�^���2�\�:���|��Lێ�B�rŵ�0�4����.�`��K�9��EV��oҝ��b9VOd>���MV+��6ճ-d��,�±������R��:pI~����O�3:C\Z�m��ʨ&�g&�x����\(��
��vu���a��er�1��Y0��)G����\�F�ǌKY�f�L���]%lS�MƄ�Ya��� ��Z��#�9�_K���<���Զy�0����s��ؙ�Q,gګ�cd:ӷ�K�I=N���U����o�B]Q�@*�����}�Zno~�AGk�h���37�&4/R|RҌ7��]�����R����qUTM���>�:^�ne�b�!=���I�i[�8���[(�8=��yi��Q��5�l�+fӐLT��|��3�hѹ���qz�������=\n�DP��B*h���1�m��K(#�Ѭ�Y��M�ӭt|	sR�|mB�d�p�4^u]{����O����.���7�H?�3��}��E�5	��dq~(��ψ�X�W���"]������63�G�0����%����h���2/���#6$�fC<��΄�FF!�h�o��p�P���Z$h|a@ ʯ�u��Ҁ�����g��_�'(��=Dpo,��ٳR!�'^�X-i{���ii�]ԈRU3�F�FE�͒�0�R��]?]F���)8A�%i%�k�%��(>�U�-�Σ=�G���L��yH������N�����HJ�auaѡֆ����|�L�_/�%(�*����[��HY�1���3yoL �o�-cٻú'�4�ބ�ON�W��V��0�<q�H�%��Vqc�p6��j��usC?��x��;1�
���p���>�����t�����:X����8�p�Ax���4�_�O�����Ƅ��LW�c��7�=�9qغ�KN Ɵrӷ�`7�ꌙy�A���57�d�>�L��sn�ԃ���.��q�F�o��v����MF���zCs�/UܧD���yM%3��[�J�V�q�`�<s�>>��#�QG�d�G�˳e��/~מ���*���e)/� 2����JW��u���#c`�yi���>�aA�1��#��_,�<�P�K$糄�{�6ue`'i�n�#Gv�Pffn	��[�f�"qV�qn�ڸF��5�{ gw~�2G�CƼ4�\DQ�dz��3�������V7�p���ɺY#��3����
g��E:������U�'"����y� �/���"-/~wfFh�L�lѽ�O�0����;�&A50eN:i�\�����l�ޡ�2��ρYB:d��O�z��P�Ǒ�	�	�p��CMӌ~L�CN��f��`/�8��O��;�ԟ��a��7P�şm�8�c*��@�[�.I���&L�GF�}�{ �]�M+4��y�y�S���b��f�!%r����7"[8��N�GBGADl��lc^��H�9�Nd|�A������jY��KR�O��KM^����%��1��i 6��\��*=�-��&�J��5��\b`]G����C\/�1��F�+�b�z��r�ͼd�̊o�X�"�ҤYDd�o��{hTzI��4�a� ���#�	�-Lk��{�k�lL�$���"Z�]K������;���ҷNS��K��X�-�i]�"�d�˒�״�Z]�x&��̫|F�Ji*�%�ȴa�/���?�x:�Ȍϱ�<���5h�:2��sPЫON���/�����Vn5�Sj�}�z�?
�����@F��A�=�D@�n���cy��@a�Tf��w�������Q'2�:��SD�G�UJN�8�[�A�������A�\D�FOR%r�����OisxoK��.:��wAr}�'����P٦C��g��=l���C�eO֩sQ�'c�֮���1�Ƽ�����$�z]�~�B�1�<�g"3)	ΐ<��/�o���.ul$�9���4���o�Va:��x){�e�����<Ƭ�W��#���rA~�_L��u9� �E�:x����"��2Ff꣏I�P�R:�Cj���)���������H_(�;Mɹp7����X�avS��Z&�Q�w��gfPl�)��`UwȾ��v\��t7M�>��J0{���w~Zlˣ��χ�w��~#3>��%-˟
lǙZ����S+w�9��9ǔwN=��Ee�yUn��dYʀ����rF�]��V�m�G�g�F�)d:�e�_�
�5�P�;�u- 2%
(���x��w�Nu}��9�p�`�AI������K��e	�Y#���s�)$I�q�9���<�|_�-�-�����6�w��.bX�[gm��9��>ai]Q32�2��b��q�4����n�C��}� /��Z�{����t>w���X��.�\S-�q20�/�wV��`s�y=I͇M��j2�9�)��IŨc�e2I-ٟ��鲄ټx&/�ވɌ'�) �_
�V:_��F����
<���[�	�o/���.�qTajvl��cP,�����JT��)l��B-ð&L̇35�d]t�cPsI?��n,J�i�SԐY��d�$�n_�����ŰG��\���e���O.jBڕ�2#��{�PІܴ���+n����,�F��������'�z�$�p������C����D�"�Trn�yvXOH��՚�����2g08��_j�Y�n���G�Y�/5��PO�M�\�K�͠�|�TO&���9i��x9\O�ŧ�f�З�]�����o���c�M�)�����B7�DY�j�%l���:P�G㡂����A.:��g��������F��y�h�\���h����m��f��:IhJM�����%��3��m�ޣk]��+������^1.{���.(7�;^W���Vc��x�r��.J�a4��NVwL���0֫s�9��y���<�߱���0ު�p���X����L���u|��1�W b��_0օ���ˍY�A���1Ȓz�O)��B���%H�&*��-Ӹ����S�<��)s��<����#}X�'f�+%� �^RM�\���y�sJ��3W��}d��)L-���a�̼n
 ����;��Rz�T�8�(�ta��l�O�7���BP)�W����ѲN�8S>��X��⑛�o3���v��]V	�&��C�rT��Py��UK�+
ֺEsn@�S[������%ʛ����o�b[ڇ�G�3C��|6��0�T[kDq`��8w�>��@hD��A�Mi`>SZXF�9Ɩ���Y)ژ�2y�HQ7�a������.��1)Ղq"�wg?�F��� ���iNf�����KY���M5])+
p�ii��fK�s#�p>�4]�$sn+	�둫O�m�{�v~qM�3�t�Ip�>���u����!j��k��P��3���Ls�Djg9�N}a>��c�M�"��?掫���B�z�TTeə�9j{]���z�����Z���*�ǫ��bg�l-ʰ��9������$U�G��O:���#��v{�ǛʬH �]�|��ί�(h<m��̸�+�y5<F�s��]�[[R�9�>�O%J�~��I�Ѽ�(a!���3L�����:�?��@Z��J*e�&F��Z���!]���`�F�;��M��t�T�9/��:�yR$Ӑaz��N��9p���8���Α.Y y�i�簍V��0\��*\��PP��2l����^럆��8\�gׁ݈˨Oh�0�_���g����k��G@IʬP�: ���������2���~8�Q��u�*]>|��:\������;>�k�ܬ����&D�H����Vͩ�b�QB���#N�r�i	��;�/!^x��NH��b�o�������(�14�x�/r�S?xqNC��	��%�E��;���c`G�6���Բ��(׋g�;c�VW�1��}�X&�Ϧ���-å�7�bePd���N�fB\@���{��w����60�-�5��v����~�|�2���w���,�G����3�D��Ae!drg�:�u��d���6i��C�)8A\�Ȼ+a<A�j˴h�15�<��/��$�`k��JǪ����Qg��Z�3֋%[��[����6�1��%��g+Eغb�:�,��&�.��H���Y��T��0P��e ǣq1S<���n��ઽ��v���h.�=��Е�p0c}����BMU#X�0�i��KP?�o��cfI�5T�I�;
�X��O)ڏ��s�wy�\�*K�H�W�!}�`�7���jl�GcZ�ӓ���Ǚ��ݴY�|V���}@����?����z��;Ǜ�ް�˭�Â�	�=�g�1&_�����(�a���-|\]_��d-��!�lp�r�؏���4���:T�������H�~�%���9��곺T�\� #$H����q���?7�����U2�m����2#����L��aPV07���\��()R�1(5jW�v�0U�b�̫�$R��J��{�@Ms)�nq&���s��Ή��K��ˍ�N:dv�v��	��%�^9F��'F�$��e�Kg��_<�)�sj�~�Á�C��^@��	5�F|��`�����|MP�\y�l0�ǿ}&k$[`������8�!Y�miP��䝪��>�КGV���D܄o�y 
��,�Z���4].^����9'ڃ������@>�Ѩ��+F�L�Q���s�.�#Y���=r��0��^QbF�W�ud]S͚0/��3�#���D�*��1� ���u>��S�s�;���l�h�$`;5��m<]��i������im��Ұ���ZL���ON�!Z��Yd�ϣg`�F)e�3%r�:�� &%��sd�ga9I_��/�Nͦĸ�7]u�P9�F:� �Cq%�T���`��)��`=��a��kC��frӟ\�2QI�і? G�T�.Ƥ4EuH�Sݬ��t����è��°�"_Z�BkK�q�HORBU�w�� �i������|`ٱ5��_[�L��
C5?{#�铃�>����Z?ύ�[�L�=q�|��9�r7׆�I�{��LU��j�	�̐:LA�JkG�.ؓ�u@X��c�K�U��ȷL)j�1�ۄ�B����I�z�t�y�����'K"i/����	k����wp�	�4���(�
��6Q����(�������b���B��6q�_�3C�M�⯰�B�nLط��hBı�����R&��bs{H��!K���aJ�̒�}�e���D�l����qn��a8�m��\�&� ���.�)>�lN��+��F빦l��;HZ_��n0��l�>��Ah���w��8k�y�����g��T�)聏�r�3jY����m�C*� �2�cٻ�-V�zj11p2�mey`k��e��}�e�\:t^������eO������r"s�3��^	�W3Z.��w���U�g�W�k^@נd�a��(��'�K�G�ctkV��XS�aσ��
n��`2^�R��ç�JFf���JgX^���S���$,��J{����9�9c&�S&s�4�Gec���"+TFa�\�:Z��] �t���MC,
�۶��Fτ��'K�1ƪ�#;n�v�-c�ےm���w;>I;u�y�W��:��a���(�����>�N%��J||��G��5,����X�d�r\,g��%�k��If[���t%
w�Y�81Gk�k"�th�j�ѵ�.������H��롭�Kd�-\[�O8���	�����i^N)�]C���ø5I�#��S��w:�ȅZm�Aι�������k<���y���ŷLKH�����B�=j\�^��� 7��o��V�;�A'�J������5DtY9i1�i0'V�O_�3�����p����Ÿ��IB˖�9��0���¨�`��
v�?�&�0�5�o�XU�Մ�:�YZn���!�� �&�E�e����P�"�6mJ��d���W�Y��6�E���$�O�_��O�k����_6��'���GIT�z�[����� ����D^��g{���>2�] `|�uZ�N���0�\�''b�0�נ�fl^��L�2a#!Δ=��bnRB�3|�0񬭂�{�1;���#A�s��1��S9qz�veT��S	w��׺f,"j�B���m`�~pw�2 S_��/��ղm�	�Y�b4Y�t�Y�Ф޴���$\6Z���t=�U0MIU�İ��1[�`>�s���ȜnہUbU�g������r���?�����
v�܆&�,S^�>;I���3�]^N�>��F�;��� �V�w�j�Gӈ-�?�d��h�B?��]0	��W��`\�״	c�E�v&aY~NY(̪'g����n��%m��dA�̈́�J[�+��5��c�F@�U�X{%i>.~W{��.�3e�K��'׬m-d�35�^-Gћ��'}剥�y�r��S�G�:����
���n��p��o����L�:K}���V�ѱ}��mH(A��i�;��3`���G^�u�7�F�ܳ�������6H߻|����AmFi�!���A�e��r�g�����B�#Ou�L?x��˗4		qVə$?(~��c�,�.��۱�S�/5��X��aӞ�ｏɋ��h�3ҹ;	��!2�h�P�:��Og������~����W3sE 2xE2�W֝�)_��6�{��zO�d7��\�oT����Z�"Hf�nw7��\��
������`�^�V-�7��ƺC��lQ����^�,�sNXoS�#�a5�N�Ё=��_�u�.اr����������g�KD�n��]��AG���
��װ�n��ۏ��*�B����d��K67�Ua��h6�1pkM"�>#�Nl~�T�Hi#�ڃ@�Aff(���1,U�L�d�g��N9}/������.2���4CB�H�;�d�{���a{�jh��-|�� hK�h@�Y�n���q�l7�(\#��P|�xj��կ��F�����Û-�yx�̺�Y����ı.�!bT脥���1�K)��Ǚ�L&��ד'O����/��EW77p�a���H�����^�:��w�T�U�h"q��"��,aa#�hDs9p�3 ʀ�>n�3t���Q��R�D�{`mٰ�#�Qt�3��.�c�Z|bR�7%����0�~����3�����{:Q��v�����)�'LKݠN����!2)�_�o��i�4���<�����Ov$G����di�P 
���&�����rnfm����?���lN���̭��p�CNS�����V��UOgƹ{DdF�{��U��	�X��Ȑ��{��z)��e����q4�H�:"9��V"A�Ũ*F��6'e���[K�v��TX�9��օ�1�X`�`
�s;A@���f�̍ɠ
��У��E���*�H�$e�Q@\K;M�]�DL}�=t:]	��$I�6�>D�lpǷRt�>J�J�^k9�~Ц��6ɲ4���|m��,	�掉�f���q�u�eX�x����x�0�}�S{|�H9�k�2!��L��i���!?���}�RxRb��� �'��Q)Wң^[&�I,H�_����@��g�ы���0%��. K���Ye�[��h�͊��I��>2�<7h�p�n����0��a����(
VJh�V���T�i�$�J�$�2q8X�X�kA���GP�|��{X����|�jΗ>xS��z���Ǫy�e�s�r�,�!iw�&I[�� [@}���u�R4pI�� 7ݏ�n=E�a��*����i��֒���E�f�J���rV�����9�n�$�(��۬���l���猄���o�~H�1����
�RQ��ݬi�e��y�p��q��IS͓�#I���ZN]0☥{�����yw֞���6U�l��i�Zݨya0gC׵�d6�^,�3im�ę���� zm���L���U~�>	�<������ϰ�I2�1�NJb�8�O�����K|2bi��hdfK��K�}���g�������[�l��C��E=�\�ʐm���KN3�����\�v-2]IDK�qT��a�vp�%^�к�x�3�/N�q��VݑREu��]���nI?����ɣ
b.Xb#J�������dD���g�e4y�� u,�D�WEb����Q�h����u��R������;���E�y�fu��/ <�O]=޺2 #���ZG���ωq��4;r�U*����b4�͔zF�Y����e��y��Q��m��w]��#oX�`{{������1���yW�r�z�x�z�����j�Y#?��9��m���J��K�j�*늃��ֿ�vB�3�����>y���j|��!�4�9��vs쓑�MC��:s��;�������T����[�18�s4�>L��M&~!���/��S�I�6(">�rMs��;�ĩ����c��#J�����fĥ��^E�#�:WYY�+Q�̗�����w�z�I�GS�ʝѸ�/���ذ�*[�q:
���	�nk��^�c>�Rsf�����X���&J�٧_�T=J���p��ő�b=Eb�}�����P_=>ID���֣���:��Iym�K�ٗdK&�U��Ì6ű�t�8A2�O.�h��ځ�V���}��������nbo9LQ�IX�`��1��3����� Z
�Z�߽
%CLK�AZ��bx�G�{&<�9����Mx����R�m��^�O [@���5�Y}s��<A=�
��za+�����cI�}�{�\A�d�l��;F�#ޒ�Ra�j6O��ݛ�޻n�<�O�T=i8k��y�^��ߑ�|����Ѫ���z�z���}��U���Y)4�wYa��C�ǅ�Vc����A���ၘ3uВ|��4��ؓ�t�C�K�^�߁Ue�D�]��aз�� L 8�!��mxLn[bAU���t�cbS1~��d�Ǻ$��r߱�;]r��4��Vq��>I��:@�\z�\�\��PO?�w�)YC�Dm��+҇�v�Eĥdn�k*�2�^,�̱�mx̎u|���ˑ�ڇy{%��ᛨ��88	bP=9���C� ��j�  ;p=������3L�)>.��Rr6Z$L�$%I�%Z[�(9#3��)��D�H+�@��\pヱ���ϧ
�\q�%�J�4!�l��UZ9֝#�@�A��^����g0x	��w![��6TT ���J��MG��>���!�AJ��0��3�\6��Tz�c��sq�&����ɇ��ѷ�,�a*\��g0����^+1>�*��/q�vJx_���61ؘ����I��Ҵ3#����5�c�a�"���W�7Y�A��r�=˯��|��υz���W�ߑ�i?�z-�Ln?X��Ck�%0/�:t���S=Ё*׶U������|� ,��7^�ah��f��ڞ1y�O�(8i�Icja�� eDhm'�x�3S6�`��L��Xk��p.ez��k+������(e01�䏅�c:�A~�烖~�8t�y���z ��i�[����[��[��_��u�����%g�&rKQQ��q�	H�Z�꟞~�0sY����P�ֿ}�`d��G������Q)��6��8��Q�f� ��Á��U\^=���Q�3p���'��	kM�(�\0��d���j��z]h����vS�� ��2��|�l�<��̮��[�>�=�v�k|� ,+6`k"͸3���Nf ����g��60�$V��"k���>-�3ѳ�Z<����M|`� "����O�s�Ä�|��>>���PQ=�)��]��(�3W?�|K��:�����[�&85ߵDC�X� ����b�f�8�	1����CQ�D|h��0��/)�8^7�3ܔ�9Bz���Z����gd +�sh ۧ���rm��3���R�$߱��0��PC�U�t�g;�U
Ec��'y���ŏ��J��S`��&,��ʹR�T�� �E�:��C�7sQ��9Rb����K&�J/FK%��A��_��,���LW
 �*�_X�2|�����ժ���/�kE������ǁX��;�\��P�0���y4�n$7܎�6�A.P/FR���'�!\]C��w坖x������D޽��l�[���b{���B4G2y��t��;*��|�h=I���g��}��,_�x���Lg�<� ���j�������;�&G�q�R� [����M2C��W<J6� @����w���d�G��x5�-�����{[���-�ս��GX�a��W�gO��ȋU�O`U�M<j��b���`�����ۇ�ϕ��pw�ٯgOf�`���*�6���s��{(}�z�d-g��"����=�������4�T+�u����~a ��6eq_\����Q���ed����}�G߾5�-bP����:�R��Je�l6�P��B���(t�%�hku8
e�d���?t�8�8�VuZF�av|��0������,8�����z^iT������*wV��0�@�"��K�I�+�|���ӦA�t���{��Q�5��A��$q�z����P�J?5d1{3��Y���|����ֽ&<?(:}���(W��QUF�\�4ܙM��N���>��G Y�\��ˋ�*U:C?/�9/_Iz��:%2|.k��1�j(p��q������SYF�~����z��(���ԭaP�&b�]���u)w�/��҃|����0�Kj���~E���>����v�p���z
�I����cT�bkc��l��E���{?ƣG95��P�4G^��Qj�M�����f�,��dɓʓ�%T+�ciK|s�|�1�v[��h#�THU�ʷ[�IO3Qf�p���e��Ij��=�?����<u�Ȉ8E���Kܨ
���ŧ|��>��|CcF�|r�o�q�h�B�\zi8�L�D�|�����[R�(����,�G��$^Vc��=����ʟA�Õ����Tԧe���է�R��Rv���.C̙�s�v�C��D7PJE�b�N ��a���34zV�U�yQ�A�v�6i�	;�����,�Kϝ�=�:� �:�zԓ�#����חU+��2)n����B��Uw���Xf�b6�El�V�W���E,��F���Q�8���9i�TF��f�2��M�
�>IL4y�!�O~����[R�� ?�Y�KS��$~��2Q���J7v�={����$5u$��T�Q�����λE��>&I���aF��� ��<��/c�d�����؃i9�2)�pUzV8����pH���d�4,����w�Q��P����2 ��:Bd���6�����ʟWI�>U?�����a%�Ϻ�Ǥ���y�Vi�p<[c����0G�Zp��q7ۈ�=Sߞ ����,�21|{��ٱ��%��f��b�|Q�A$s����c��&�3b�`ϻJ(E�4X�	�b|pXM(Q�	T�y������/m	N����γ�X�'i`�ܺp�# f��Hn�Ą��u6���:��gehQ���M�2���h�Z�<`����J���U{Hk֧��0�F��͒���d�.��%!۠ߜ�T .⻥���-���!}��5d��$�qA�B[�%0����Jjo3%�$�^����]�4A�QW�R"!և��8_0<c���Q�AL���{9��j!�(4�a�8r �'?ǳ�����fdN.�����KL�>�$�SG�ܕ�H��P|� YV�
�k�����y���8��4����7;\�\�I�m�<L��'t���S��І���G�v�-8q�oVY� �&ޜN�sD�`G	^3�!ޟ[�[;��v��ѩ�5����@� ��\ް����3o����fd�{� +��)`777��a��fo۾\�r�<p��y�;w��X�+��8&sX(��g`�QnmmɫD��>9vrI��N-f�3 �S.�:���}������"y+Q�s�5���X���䧆!2�a�H_�,�R�<S9�ٕC�m���Ic`�k6J�	aF�2�����\�U�v{�ޅ�U!Z�Q}_�X���KRI�����m�����!*D��a)˙�3���!s�N��m��n7i�Ӊ=	��~ K�� �O��Y�ǰ�� Urz
�:�0L.�����v��r��׋K�pнxgj�<�|�Y�.]+�a��l��4��g��)G����F�tz��Ҩ'��4{���7v64��%0L�����T��! ݸ�ٷ�ge�r�!!�c@C�|/�8%<ܑqʥR�Ji�5�6�@��w��y������Y����-�;N���z�ĝL%hw���X--15�YXX
�}���o�a�ԇYO�����ah��4U��Vʪ�a�Ĕ������":s v�f~CFr9+���c�]nP�J�E�)�y���W�����_��c��5���X���+P֬�X�[��T�}�B��,�Ġ����,'��fe�rN�|���gf��F$��n8�R�c7�2)�سs�?�r��bο�D�ζa�z�d���b���s�av�ᠥ�	'j�uG`�c������=C�imR�g9��� �q�/T��5�vzX�?p�x��"I\	s���,�2��|���fug�J���T�2E�,ѩ)�����s�0PAfR/�)�����C�9�s{[�^�e_+�=+v�k�i�r����"�I�:^�:�\ԩh���PZ��N�6Զ��ߴ����/��Y�C���d���}{���/k�=���ξ�.�	����;�J�}���rjB�`9��pǽL"��e��sǹ�(��������2 Y�{9?� ��gƪc��pcH����@��T�u|p��'-�����A��7O�,�+�?�B33��0��~-*��tJK��Kg��[򍜁���RFT���|k�������W��޽� ;0s�`�oÜbDƴ�}v��Ȝ�K���w&�k��r3�myF*��b��oGƐ$�P) �Nˬ5`c�$�C�s1+�	���YY'��:�l�<+O[!x��t�i�*�2���K�g���B�opA# f6� �u���6�e��G��Oy��;|���3�r$Y=�E91�)�k�1� K�ĦA��"�w<Egԥ�4� �3"����M�7\d}��,`�x�I`��E{�v1�)����T�Ϭ��?�"�y�ӌQ��a�.�>(���2ʓt*�=�����~�	32ވl��au~�6�t�f7��Jm(�ؿ�7����S���[�ަ�������4?9�ˤiT��=s9#���|h��|W��F%^�3�WNX���qI�6��E���)����S]�����MF�!F�<˘��b��Y��ުKzƀ���ŶNq	�K�ӣ$J�*��|X{R���t��><�Wx��GI&�Oe�ߌ�k�@ڝ黬�CT.��X����
3�a�,���}�=B���l��wMfu�>>�gȝ*�]�]YIdy�L�H\��{T��ѰZ��.!�.�W�c���7��c��k�ö��'�����G� �� p(rWL���ٌ�3p`���H���T�:�AA.��ռ�|�C<zA,�؆DDxe����t�:1p�d��w��=@_���ח���U��Q֓x7>����.�:�����a�����sQ��;�ɳQ���!�i��[ꏳ}�G�׆�hO{�?��B#۴C��:����mX��H�2�پz�h�g��}�N� �~Ү�*|c�P��~��W���'�}w�0�ڎ������pT�oD�	�5g��˨h���ݽ�+G�1xΝ
/u9>��<O\e�8��B�3�=�JF/%�f~�Fk���Z	��*��I�ZG��ט�z�o�cX*����F�� ��u*�Eg鏿n�Pt�/A�����۳�d?��~�3�߂��?�ՠ3�`b3נz֯a�Rr��zr�~���g��:,�}���`��z�J���Z�0�ϹM�
�M�ŅB���p:�{��e�y��@^�{��a	�	�c�����d*�&V�� z �S�s}F
^Y��~bVc�8:U|V���y �C���@iIx�A9��;e LF�ie�Ѕ�5�� �؞!�B��1J�X�43ȃӰǻ9������C���jV/K@Y�����_�\��3d���t�y`�}��(M�P��CWC�J1z�m��h��S�c���92�yR7JuvԤo�4�V�:�a
`��*&A�8/��;s˝u�p(|f�L�P=�,���� ���G���Y=GS�_�(ke s=lj�c��s.zM�������52@�� �� �b"�g+�.)'�Zi%�$)$$���y9�����#8)㥆�/Ke˗��@��l��/�IX���	n�Og.|ܐ��5��G}��P�v�w6�Ȟ��~ߑP�R�`���{{��{��k.f����#`n����t��Tu�{14g�����S�C��+Î�����1>O����h����$�N�4�1���r�G�⼾�{�z�{��z�����Is#��/�S���`��� %�`�Ƈ e䏼�DkK�W��;*����SOqN��5�Y>DTF)�!S���!�X�Q2I�_�p��֩�挛t�]�ad�(�3 2�S٦�ψtB�9��\��U�~pQ���k��ݝSU?#}���2мJ`R������@	lO Vz@{#qp���)4@��p��������
����.n�rZ��Ҽ�=��A�~�]ޭ�[��`װ��:���=r	�Ym�
/���;:�����Aʈ 6���lk���ۑ�IG������V]A����B���f;��V�
�p��^���;����:�
�o^�չ?��d�����	�P��ws�h�k��A���[��9%Od��� ��N�I@��Bǂ�q�w�t���^׀xb�6˥
:u#b�Ȇ���yMT,�o��A�RP���u��MT�5�E���V
��\�8�C�2�"����$e���^�V�z��g�H!=T�i���T��0G�g��W�4�I�*�1���X FQ�S'u����vvvM�q9�|#�\����h��&mI.�pn<��j.:B:ԧ���t�q}�V�eڝ.0<�d�3c��n�m�ns������ڜ�&J�q:d��;�`�rv��1�T��s�赺�hr�m��]OL�z�?E�G�0K���9pt$0kJ��{�Al�[�>5�sr�������|�bmm�G�����IY<�F���0z<̼��d�xㄎ���V	�h
�2(��,c�`;u[��Gu��1�l)�c������1�'%�c�rP�B�;t4��p`���q��=�YtV[�qjm�\�=��Ebh1��q)�cƙ�����>�Ϭ�A\6Q��#
f��bQk�&4��9�N�r��S�}TeS2���3�g##m�+ŵJ	B�Z����S�Zy���ӣ$��PðqDGC��H-"�*���p�myV�^�3Z� ��2��zJ]�_`.���̞�L\Ϯ"��D�F.	=��# �F�ٰ�	`�s�Jb72���e���S+��.�yv�qJ�LBC0c��aZC�-��84��0�͝q��#�r�Dc�A����>Q���X�S������0�m��	��HI[�
���*31݄����*+L<�h����]1��"�|n�����L|�:���Q�v�̧0+�H�`,��27
�����J$�t;��L��	4\d:H�JI���isS#��`kk[֌s���G�xA�(+���#�I���%ͽ	����@�&�9�% ,��L��i�%&,�#�'th��3r�|s�f�]�����d�:d�������L���/�%6S[���F��:{�3U�r�L�RMm����L��y_�L�泧+9�9 ̅����aP����/�����]O�j�'}�0#i��s3�0;3�G�F�X��W
*D�O6�&d���c�^䞍�D*���a7,�r��89� ����c�#�$ξ�
��駟���tc��k�����߹�<�krvǏ� n��;w�`��k�D�N��¹s���ǫk�}�6I&m_\��3gp���|pMA'�k�s���i�gskK,�®�X����'199���u��~��0�p��E�7�:����&�'�q������' �Ɣǒp�>>�S˧0;7#�ŭ�ױ���cs���ǫ�q��=�d���8}�|�9 ���Ѥ�.,Ù�g���/���h6(�T��b~~g�,K_=|��w�V���˗��nߺ�4��ID8$�J+kL`�?=3���i�J�"�ݿ���-���H-kjh��c8~�8gg�i4���������A�A�Im�m�)�¨����8q��n�n�ƣ�GҶ�N}'�>~�$���*B$*i��%���"�-׵��1Z�7P	�8Akd}}�H�����07��_����.>������B�lA�ӵk�hM����4V�q'F��?w�<�,��y���*�����߿�����wƦf�8omm��tw���J��3�w�H���6u*`��%s��W���?G>1��H9be�z�"�F.�_NמC&g�Vm�N9��=s��$�]��-\�0z1V�E�W��ByVϓ����3@c�a���Ξ��S��h4v����"�D�qǢ�ȸ$1�����3������__'~ǨuX�	B+�)9���w�:�ݤ��Φ����N��ɋ8����?��R�@�3)�]�!�;�1z�Ƈ���g��,��w�`\��0)��|,͞ĸ����F��C�W����y�Lq�|��*h&�i���8�� ��!�d����_"� yo���n��b�͟�:�[����&�8NN�ę�%�q����C��+k�Z$Elu%p�8=wy�7B�_$I@�e�%�n��K��	�f��SJw��#⼅ũy|�ŷ�����6wHJh+"�%�jY\���Xm����˯c��c�v�,-.	6�[�I6�1ip�d�8<�@Ui>+��Y�����47�����cǖp����x���*��._�������-�q*�,��������K�K��T1�:f&g	�g�ŗ_�s?��:�;�Gl��1K�>U��&1Q�.���ԉ�x�����G���5��Jq��1��^~������p��?��)Z#��q�{s3��w����S_WD�"�g��h���so�ebv�wp��y��ML�c��*I�c���$��o��-4��>v��/ն����ӎd��7�>2��<H�5�bW[ow��<�<�L��ŉQ�gV�LX2(2j�(/|���l'�����ԍ�E�[�ݐ�y) cT&=�7o�2�����c,�(�I��NCk:7�04Rr�����5,�>���<>��(b�4�]�$Iu�)J�I�s�>G�0!��J�8LI�BD=�&.�[`A��h�B@����z����`�.fONc���d�i�����u���q�`���눉�?��� ��$RL�o䳇ڭ�[$Y��%��ݦ6���P�d��=K�Cu.��4��J_|�)I-���f}c��5 `Fj&2d�Nmj�	��h�??;��ܾͯ����l��e,�_���zl�I�z@OB��܉%֗��3��حĆ=���F����&����**��|;��Xmnb��UYI�H��u,����^�����u��.�K`�MLK;�S�ޡM�)�H�N T��"I�C� �	"�M�%�0�]lX-��������v��B�S��F�^_�ti���G��1M�ƌN������n�`{e����u��Z3˳�/иV����;C�>U�ƺvm�.I�/^y�X�����˘�9<N�s���-Z�ը���q��x�$���$�PӜ/3����ښhƈ`�#�9:�|�[���ZA�;k����ll�����6�wש�m��е���|K$����a�$�-_>�s��� �2�:���;���$�ϐ�]S	���dϷ���Z���	S�1r�i�y51�p�>�6N��Ӑ��ڸ3,ASpJ�}�)�e�v��Ia9�Ƣ��C&�O��KF�[�G��-�����~b�֓J�GQ�A�Q��qr�;��ŴF76Vq����ͽL�OQ	+�"�-��C��S�A*b��&q�gp��4oWM��z�՘9K��7ub���6n�<`�6��k�p���m�����a3�6�U���1=M�hm�������Hܸv�'?=	K���,p�ы�����!V�!�����C�v�(�#��I[6e(�!I-]Li�T��|�<n|x�h�;�X8����L�	6=k�Z�q
0MR�l�����"]���_�D��`�#�
��9�&I�PN8yg	W7�03C}����<:4�[QW��+0z���Jgjg��i�T�������?����tI
��6�9��%��ˆQ(u�m�!��k��k���%��E�� pLLH.�g�\k�b�։�a�����X~����Y%ǯ�gQ�fqD FR�Xe���E������b=P��x�����U�:}�z��(w�4'cx���.�g�X���S�Ʋ]�x\B���jy���ZP���c���g���n���F,�t�&?�qf5)���(	��m˘MNO��s�ٻ��W^}�]��=z*���+wP�U��9�u�N���_��g����{4I]̌��$f����E-zo�HG�휻�{^{a����`r.�K�y�Q+�g��B	w�����29��'�9 ˈ@ƙZBA�HY�b�ˊ
�Q76QX<O��_�r
���9j�']}5����/�9{PΑ�ه��1ԓ2GP�A�����}��MB�\���j�1ܹ{�l� SwqĀ0�jb���&�ܺ�7�x��!Fs��MƢ�JM�ݺ����'����7"w��µ�w1��(��:I�ѶX*���DP������v	D��ssg�+��O`ksM�b"Ц�F����1z�wi��Ф6���]jWG�f$j+>wR���"�K�o?|�{w!,�Q#	n��:q�rSĨ��ľr�6h�X�!��+�^cԶ��cB,�p[��^&>�Z]�Q>����*�v	Ğ;�,c�s�akK��d+Je�]���k�����z��0���(�F�+č��M�-��e��'�1?='�e@Z���N���v�a�b��FWy"mLיp��c���w��S��b��3C�(Ϛ&�-"�H�^8A�I��Khx��/6zL�bвKt������XY_��K/`jz��I p����u9Q������аd$�13��h�-{���e/j��j4���E����%��Ȅ��@�Zz��L}�@�$t�AX^>����h�����岬VGNON������1mi��s��0*������Z��sPe���fO�h ��Ov���ƸҎ�Pߪ��'� ���cĤ�P��.�t���qe\�����)ier�/��9��٩�I9��ڤN����8�vWu�Q+8	� ����px���!eT�!'٩���?�jy��ԃ#�׈��'M�-���@>�b��7�≓��[����߄���Y3�#h�Є��MD��=������[r���a�RbWw��bԈwH�������k�����x������c���w���CD���H�w�-@F�4	�T�D���-��W�<��ZX���$n4,x�{'*�x���Y�RB�o���g_}�׈8N�&���W�e� ���cl���x�=����x���q��촶�{$���T����43�V��m���=���|�$"p0&��BR��[ʝ�6���_��i��?�9v67P+h�i|��ǉV��`�M�\��GD`�����B�4����Gc��	LOL���j���0By|S^�Kg05>��Օs����wx�����p��!Y�-įD���H,C��8��38s�<ʵ1�^�P)���2��{���m�nn޾�$�jb�L�����9>��D�1�Ǯ����kb$�u4h��~�m�iN�*13T�K�$i��2I8���*�`莀�.���}/?�N�l�W#��>���M�=�N�A��I$�d����}����VO�w���4o��}W�~�.}���
vH*�E�g�G�"�c׍K�����ki��������|[,4Y�}@q��}j3�+wV���99�y�IԚd��nTc�(��@X���2s^#F�^�a��g^��[;�hno��
%Ƨ,ֱ���ʎ ,�pa]Z��hC���y����<������K�!�X��X7}��'���᫻7�#�hE�.�:����`�4��z��|>��kp=���x��GVF�� ���R���i��|�@D\t���Gwb��#1�~p�,�0t�ZL�{�mc3o���_IMa?���A�n�~��*�U笚��-��\�WW���W���i����*�Y�Ư~�+쬮�y�#Q���KЁ�KD2T%tI���ZG{s��_?�w��c�>���r	DJ��j�_���O��?,6N���p��;Ty����q�FŪħ��$������&��k����$z�Ӽ�x2��Pt�D�����C��W�[�k��?��ư���H l.��&�kᗷ������
����������@p��Ck�D%�[c��&I��~�3�$�L3��o���Gč�W� ���rS��՞�������-��4�JU�Q���?�9:%�R��TG�����B�f)!�֋p��[x��}h�0jO�3��b*�|��7.�H�#���v�W��������׮���X��֪M�=��ύOc������ߠz,m���6n��?7��D	m>�uU!�m�|Ѩዯ���?���3�!]���mjk��V�a[�_�I\!�����i�"��4������Wps�]�����+�O>��mC�llc�����>�xW�1J�����b3��u��S?mo�E���aʴ����ї����F���,nuh�+LT'q��Y|��7����|���YM�C���w�?�������.Ia�L%�\���� 1j9���&���P�{������� S�1T�F�35X�j8�����"��w�	���n�Bg%�|�DzgP�&���!�g�����>�����(��^�8,�Cޟ�_6�%�W��,���ɔ�z
@<(�۠z���W�k_>譖��@�lHkvq�8^:��-.!�q��]|z�"<dL4���]v�iH��oi�8����	v��׿��?��;ۨO�шM�C����m�V��3x��8O��4m�6Ie�n\�/7�ݳ�lH4L��针'�zX�g.���2jDx޹��n~�;kw��٠��&�������8�x�����}�.>��3�����
Jb mG�2A����%\:y�'�Y���7�⋛���/	c��q%�H��Ѐ�B}
N�ƅ3g1C����*nܹ���&y�Z:���R�BR`c$����{��������z�����['�l�k/6t�G1F�??1����3�'������w�5�k�H��kFKu6陽F��3x���8G�u�ڸK��m��{W�U!��859��!֌�uz�����*�������n��8L��H4�E�`ɶN}��5����N_��<+gl_��
_��
���A���*�b�Of]���Z����p��s�:v���_�����_c�$U]#����N�-���V��/�xМO�\������p��5ZQ�0-��ףv�����I�O]�sg.a�Ē��ݢ9�Ns��ÛH�J,2U�d�ʈ�c��J���'N����X8~�$��|�{|v�6�9�d��vڢjMR�����(�<eℰ_!?'����~�������%�듘�@S�y0�O��_����q,�<���'����*�y�c�����S��9X�gj������w/����*4a+�9a�	1QU����?���hv�����^w�D�$��n=ZF�_�>�H�F�g`}GWϡ��eC��d�'�'�t��������=�*�����	��oZ��^y	o�[<��r]T2��{���?�o����m��nЌ1K�������������x_9w�������'�j�p���9���~�/���s����%"p'���$�����f��G��q~�,��?©cg0�*�6I&Ǘ��+/���>Ŀ���x�^'0�7�ı~��w��+���ܱ4Bȫ�_�D�����n�]#.�-��w���OM�/��!^y�5�Y,�t6vp��g����>�>���p�=ѱ��i���e������S1=6!z��]������4~��I*z(���-��Y�x���������YT9

؋'������O��|�;a���V�	ز������˧�#&�I.Sr��ui��᧿�%Z_~@@�qB��y��)��?��Ͽ�IN��j�拯�=b���/���MԪe9���N>Oz��e��k��K�xLDإ~_Z^��~����?~���:�FQIWt��/⇯� �fN�ض	8^8��;�/�ǿ�����w�1,��꺂�����e5o���i�����$���_��޹MR|C��0+�Fgi����wH:yI"M��V�tq��Y���_�W_�G`}W�%�\����y�����7�=����4kP/]������{>�/n|�V{K$���-���,����F��P�a�����"�\�����o�d���F�q��3�*ݥY�q�� &nfjo?�~��;8>FL1\�P�:?a	9f�����>7�&�����?����;�E�Qֈ�q���)�k'����ko�q+!�s�܉�=�A�j"�뗏��_�����U<x�#��v�V�W������x�6�g_B�}���f��:�0-G��	�߻�������b+��J<���7���� ���X~�L.`��$ƃ*q�[�z�.�DM'j��w�ܽ�t	��)������xe���	���ߣ�:��绸�jx� .�-�Go��W��#)��`�6�8�7=7%Q:Vw7�%�آ�L}y������8lY2:4�M� ��P�>���/~���_����5F�*�ƈӽ�*��ڹ0��d�����JU,��?�2�qw��a��#j����<���{�x��8Eč���$)��k$��ѡ�o?��[�io��{	Nҵo���[<->r;��to��S8>3�5��{�Iy�$�N��.�i�G���H��Bb�i�PL���"�yb�<zt�[�I�0���_o\~� �XZX"᪃m�Ҫ$��%f�Ǝ�;X�p�z��l��������KW0����A���g��NLc� fk�>>|�)��r��k�<I3Mk�ʩ�DlKX[Y�*{�5�N���wТ��B$���ǌ�_=|�5"��n�-�h�g��&�� �]�o?�?��ޕH����<�����W�q!�rkG��IP�y�"�z�@����6Iʤ���~g	���y����R�6w%��"���b�&�x�l�u�1���
����������ǡ��F�O،ժ4�-�7ޒ���霵�4^[M�;&��Mg0�@�������K/�����
&+��v[Ƙ�b
G<���{W^×7��{�o��|����'�����F��uq��'�P倻�u��R�O���	伀-O�.���v{��M�O�y���>aً�?h=��}�T9��|��8��@�m*����2�oGhE]��A$�p��y|�xW��jcC p�8�׈C=C`�]�B�@���,6[h$m"�U\"I饳����]��D�ju\>u��8]�Ak�C\mQ�N�m����9�2���1�vP[@D%���<��x=�q��]��tM�$��S��|�y|z�K��yL�
�7�����It�[�$b'}�d��$)�����%<��"�𞜘��/bI�Ѻ�Ձp�M�@R� �pq�4�/��֍OEjC;Ƌ�/�U�Y���6�l��IZ���"Z��Ǜ$�|~��t�Bhf��^:q���[��q���m�bl�~?y/�_���wŷ( ������˯�,q����ٜ��Ǐ�165���_��D��nl��D���||	�\�L}/c��}�5K�]Y�F�S5�x���&V�l�bK!^���������k���ْ��^�����$����_�HL�9b�%�+�P"i`}s� �+ľ�����^'�|���ׯK�,��l���� ����M��F���[X2��������Nae�!�n����gC��b4���[DW�̏ƞ��B,�")r�X�nl	a��8^>}����Hk~c]�#�D�%Z�e�<I��n�\}p�qG��/Ӽ������"F�� �HId�ɹI�q�1�����Ƀ��0�)����ʥ�Iw��:`���'N���S'�*'F}�k�@_h���jɞA.֦�����5���Qq�(qV"0��U��4u����(��A!7����!�yfF�����!_��s��]��n��d�,��r��r4Hqw����Ԁ��z�/G�'�NhC�ʢ�D)*�q*6�;�7���������� kϷ_��T�	l
1��C��g�1]�D�Q��.Ѵ�������=^�ɱ	�>F\�8ڴ��]>7�`��q�i�<z� 3�	��U�Hr���!�I���c'�@�9�rHqi3c�Э��5��E&���H�u��{��l^ݣƳjfza���1"�t��xUz�i���.ƣ)�"�ca��o����N�X:�����A�8�2��/�?��s�s��;}�>x�%6�;�'�3��ɳP�����019������D	�%i���%|��'�Ys��'Na����31u�6(�1���1]���J�ҟ!	�41�u��{�P%��W*(�e��7�P�)��y|7Z�c�/Ig��E�Y�H"�L��x]&�4��'�q��)T|EDy���H zr��e�<|���iZeqnѳ��S8I`tz�8޿��L�Dt��s"�m<&	�����������X�M.�ҹ�ޥ�U�B�lsnvV\�6���TK59ڥ�a���1,L�sS�N�!Asf�a~�����$�p��9H��h�Aknl����'�51U�m�;�N�Ǩ�c9n�k@f<���j���$X���,nݼ&`�gng��S�t����qG�h4w�*1f�f�9���ctI�g���pbnA��vIb���&jݤuR�Ǳ�i������K��6��_�3�8�&���{�����"��)b���ڦ} 
C��g��L�2Y�{/�9mpH�ʝ�;��S�~U�����c�IT��%��M��p��;�7+�!���2qS3�U8ph�R�G��)����1�g4�~�Q�������Ny��6��}c��w�z|���Y�hk�
��<�ۣ�!$�-���_Z�01|�z\���k�F>� `b��"&�TQ����ؘ�x�Z��
*%v�-�߇lV^�e�@�8c�$L�gE��L��ŉt���`���힜]���A��h�R7&�|�E�{�@�A)B�1��c��%N;�s�T! �;�`���6�z�6z�r��	d��]��R��i$�f(!�VV	x{󘞞!�+s���}3�c$����&�:8��D��4IVcL��˚a#�j�U�&I
<�����N�Ha_�z�F9pc ��*hu	W� R'"%n8���a���s(&oq�Q%z�$�wmSv��P�+AI���$lm�`faԦ��bc�Z/�h�ƌUa�l�p��D�zV�N��MH�=1�3�2�ή���ؘ�����
Ѻ��i!��DN�(-11;��Z�q��n�J(�U+P�Z�d�	T˽
��m"�46�1��4IZ$�m�m`b|�A5b�$�I7���2�HڋX*c�7[>�E��3F�]�6I<D�>a�6#>T'1"ɫʹ�z�����3��Ǝ��ƾp��N�&��qZ��K��غ��B@�Y��T�qۉ3FS}V�Ns�_:=�
1;9��Ҹ���9�q�Fz��XoM����qY�^��2*�	�b���c�9렜'�Y�MH�6Gc���� 0������tyOe9��t���%����I�J���c.Ԑ�ҷ�AJjb.l��lL�8M(��R6v!IF�,*D.2��%x��!G�X�N��
W�� ���AGIe���,II�sNIa����(���	��qX�ئ]q��Ħ�0�	?��TC��J����O#�r��b f#�)H`b1O�c�u�3	v���v��&4��Ǣ�j�TXK����0HS�H|;�����`�^��)�$
MRX�6�%tQ�	P+�z�,A��H<l�~v�����q�F��z،��1)���f�,�X��Ǚ�}H�0z.�Gұ�2�V�����>\�}�m�:11Ă�E);�K
�RhNWH`"ͻ�㒕� ����$���#z�Sx�T��( �¾b<�,�w9q��L#>G��&�^9��0=���spbΗ�.�����Fl @�|���m��$��W�}�˚g�D�;�S-�t8��ۦ�DmLZ�+�k���ڭ�akmE���O�fH<M ��R��ր��:���d��I]�BN`R��� m<9"����]�т�t*�I�Q�����E��e�̃�+l.ϩ�l��D�SIh�w��v����?a�@��N- ǀ$�;,s�m���&ʑMj� ����0�͐t���m�k�Ư��Y�(��8�2!����KtG��6;&�*�� B�K¬y��܀*�
�'����F&�g|l���-ײ5��P���g&�Yߐ�#�n�%F����0��}tyˤ����$V�I߈��j�����5�/�y���ڸ��0�98-�^6i�kL8!%���a ��qd��6������8�K�&2DngwW��U���b�1.�8�*
dL����H�*�����AҤl!i� ���h>B6L�8a4��^]b8-KL�ŋ5&�.c�m���$�*1Bݝ�X�1ȱ�c���*�=J�	�D�� *s����c��^�Dª�F�5��u���>A[�|flofR��*ua2�_��81f�b���Ql"{�1g��ڦ�+̬LNL`k��2S����&�ѫ�d-�XDLk<�gu-h�� ��T�c���؂��P�8�q"��a@R�JL�-��(Qvu�T/�����G�|g�&�&��a�a�#jT"�I`���t��ŏ�H��"�xg;ݎ��0ٯ"z�2�"۟�e�rT�*�0���Oq���� ,Ȟ��Q.�.��&��C�0��}�l�c���&�cd�V�(�Zߜ��C��	u�̄�jrE�����,+*m�LJޯj"����_�q�s�D��h������{�t�`� �Z�Jd�R�F��
ن��������ښ>?Nc�K�sl��D��Ԧ����|�pOr��j+�M"t!�l8!! �P���*����BpJ���*��� ����	����C��r�V�q/��Ш��8��$-�䌎�y����3��)L���JT����$��9c+���NK$�	���d��Xo�t�z�s���L�:Y�e���$Q]z�|FB ��"ݲ
�ǆ�:>F���%�����Kv��}����ѣ5�o��\,_D�ƿof�e�][�����m��b:\��Z��0m�s�EA2�S?]_�Gp{c��m��e�elf��X�Ÿm�I��F�@��icu����ɓ�(�؁���}O�̥�IImZ_�V��woc��#��D��lp_Iw�ҨM��s�����:UH�Pi��@g��XeN������'���^����ۑ�/��+q)����ؕ�&��\��׿�*p������WY��a��0?��_��Z�]��_�_0B=�����\�j��E-��������S$h��s����b{�Sh��2�=>älN6=�e8�M�h�l��#�_�tIޗ8C�lZ�;�1�`��h4� 2�h��@��vc����$I�>�
e%V+������n��!��ǌ�s�8�p`S���ɢ\��7L���M�^6/Lh�4ΤS��y&o��s�@P��j��x~*̮�WN�be�Ĩ"��L�l����3&~"RP1`����/�*����eTe)���0��C����V�1CtD��E��T,�m�XI�8��D+��4���$�r�*��c�kF�iV��ڱ^�:J�^�uU��ğ�D�H�Y{�H�6+Kd>���IJ\�S�Z$#��,Rp�Ǐc>��qI���<90Q&[�Vז��D���0=-�&���ƕ�c�q�6���Gƀ�T/���	:�y΂���D �|ǽ�l*f�8�/�$V'h�°s?��*I��xܹ��ź�f����n��s8;{\T���*+� )��Uگ���?��ĢR��Ҫ=#�3}��6I��F�����ū˗1�́�˗��V��-v<�n৿�5��~��� �ܱ��=I�!��/>)t�䒥!O}.�c��w={�%�
Ż��z���5��B��1_����>�z��]����Ge��Y<.��)�ߠ��*-�~{���_�j�	p����;��tp�I�~�gg@���ZQ����g�N��N�B�Zg���H�rӕu�lVQձ4� ����o�ؘ��b��*�!ْ.Ӹk�QA���ZH�g�+ �2�!Pb��#�O���g Ӗ�$6K��71��b��#+:�M�,��x�\�=|��A�BC�{�8�`i��mTG2�%"$b+g?,��$1�vcn�R�R$jÈ��r�&vM���%�I∴��8b���8��|0Ne���q�g���t:��U2�?6"�y��<]�җXX����Z��
�Y�Ef����n�(JF��H,�����1��O��A��KUb�D�Le����:�ly��J���Wq��)�;�I�l�Ė�rN�H����D4������{���
S����9�\iTj6ȸ����Tz^Z\�|u��g�� ���@��z�%�����ae{-� K��Hz�2L٨��+OZˡ�N��xw���/o���'�yڽσgQ�p��I�`PV�e��&��#�?ÿ/K��JI9`.�(�*W��#_O:����-bX���_��YR�Se�p	,%(r�i��N���+��K�e1X�'�3�%��P;�XYK<?ǉ�z)�*�4B���?V�+6R��5�2.ޯ2&�,� +򋫯�ۆ,�3���
̉k�.hg����Fޗ����?�J�?"�k��~���<��c��Ld{��1��@~� �̒1�ցJ�'2F��6?Y�/{�2~O��4��IU#�]�}�a%�k3]���U�ԍ��n@l�w�����Y:/��T�v0�tX�sڪM,[a�t Q���(�}-H��CY�.�Im�J�rfک�8��i��U�v$�7��!�J���'�����~�-�9T�'��~63.��������+[�Qk�ZŴ-���˱t����u�F����N_q]��#�8\������/�����%n>��v9FS�DT��!ʪ!_�`�}���ֽW����v|���)n����<����������&��Wæ�S�'�{���(���"��x�p�PO~L�ڭ�`�T�R$H�g���s�r���g��>C��.�>;�Vbp	�dj2.G|tqN
���}qT.?��#��)��+�W����ɠ���{k>�gh_ұ6.�&�Q��p�.EF�U��l=dU~Ϥ���c����20�}	�X� 뇲�^���P���7����}�d�J]y�0eBa鬍���3����ef���h��{���������'qݒ���_v]BgօPi��E�H��Y6���C���c�\��O3���YYdVK�θ���C��o����^��"N��Ԓ6��
���:>��5���#\�{e,z�<f����:A	�̗_�ZIt�$?�m�www�PM|�qCY��*��D�n`um�ݸ��i�dm�O(I�$i^Jݔ�)�܆֖��K�P0_r<E��`Z�@�%�v�.\������^=vS�3���i�/=�Bך�N���[f��|I)}�U��N��Q�����b=b���u�R���]&pg���>�\���T��OqAV���c�,:v��%�B�a9Nm� �y�ٲ֞t��6��q�9�����:u��q;��b;R��Jq�ͳkfo�/'�T	�&a���8�ztB�m%co�$�]c#�ٱ�]��3%�6J���N+`E2+,əWK�����`�E��Z��^��<n��Ȏc����@J,��X*%��YI��J;5��*������P�8�i9qL���L��~������&��h]�[6����;���<v�S��������� �zdYg���2/
�N�5\�$h�6�v���{�W��㻸x�s��%)[�>�Zõ{�pk�d��IzӁΤ}�W�E^�!�Y舳���J��齏�۵�{~nGh�[b��uu+�mx""���I�� ?C�I��ʧD���s ��vK�H,}U"���M������}�������t�aL�������
��t 2����ԉv�f:%s�%\}E�wy�3����S�ˬ����L�t���Xz�I�6�&O?F /��L8#7r�㘉T`��kw�y�(̆�!S�5"�"�0_�;���h���4����FbȞ�� �.�c��!�M��
$������6 [#+�ضX�#��$���(�\����s��@�a�T�N�ܘ�3��J ,� �/f��� XJ��Z��b�`AJe;F�É	wĿ%�*ځ�ar��2IO!���*mu9@-[n�b'� ��rB��>$f|Tk֦[[����I�xg����la����X��U��)s�;�W��%�YVJvH ���N׻�f�R���Z)ֈ�誮�%b�I����}�>&k�2�w� �a
�8w_/�c�h��A[·��lg����8�P�!�\�v���Xk��<�P������:�L��MP:GpY5�O,�A$9d�/wV1Ȇ^�(��Δ��!�n-,��=�nLoS���g@���,A��V��8UAx��K"���|=)k�n��V�C!�������z��H�����ȡ��[>bIc����д3I�=@kZY�6h��ɿ�^�1hH�@@;(0i)���c�O��I~-�N�����:�ͪ]���7g@���a��и
t9	�m;?�j�IJ�#���uD֛�B	t q"�nh�#ފ-${�n��ᒈ�(ņ��=�%��y=	�e�̵S R�G�o}ߊ��IS �ƣ���V��,�-KfA*��d���$�f�������1v0Fz�bY����Q�9��Ѐ��Ҕ�G�0烰���Ge}��&����&Q��N(����grnF��%u�� @��;ⱻp�;��L{��80iM�SY;��%h���`�f\�>��<����\q;;�6?2m�r�7��T�����2�F��Y���@�q5w� 4�G�G�$5J�;)�b+z��>�W��lsɆ`L��\؆�6��6���y���A�{�߯��'�n�����+����=*猳S�^=�A�'x��am�I�'{R���@a��Q��S#�__̙l#&�e����shG�-Aa M0@F�N�p,��_ȑ,�Z�,�5Tg�S�=����%�	KT(��q���O�j��c�lI��'z�/Ie��U@h�T�v�%Nہ Y��qO��c���Y�8��')(o��ؙ?�'"��'��R�H��&|��&��HrI%��r"'r2�R�=�ͨ[ʌYς�(0��B��ʥ����\�5�l>63�HJ�	weU���=��C"[HO#;wJ"ͫ��p��кĂ �qd��ӆ1	1D�z��K���@�� �gq[#H�A�8�wW��vRf�Qd�dtlZ/���R��5�d})3`�[<Ÿ��Ҭ���_,����[f-=�����Ӧ׭:�j�"ktf\��9�	e��f$���.��K(�T��\�ܶ�dzo�Swt)3*��AEg�tt:%�:�J7]�'��}������ܻ������5��9�,��@"}��J}D� 浩x&8hd�������Mi�<L
�U^[2����^�ґ8 �?N�α�x�p|�:���N��&�OfR�î�$y��P8}>�N�J��IW�	���L��Db�qx",��YIH��,*7"�U�A�3o�#~����!�Y��H"5�I��]�׆}�r]s�.!J�+��A��b=���#�:a������I���tF\�S]��<����|�})`��d�V�T�%;d�t��_��4���%5�xl�A�P�,����y�mÆ9@��86|�Pc>&��,�bk����jS#�)�z8�:�/��4�<�"��II"0R�=���%Y��ٚ8�*�����F� �!��ƃCJ��6�Ĕ<3pҋ2<Ce��c�P�&V�v@X����FN�i�*Կ���,�?�j����ʭ;X�߱�� *�64�a�*e�v.��El�$c3G�u�3��sZ&3�?{od�u�	�̷�^�¾��}�E")R�.���y����{<1���D���#��vL���v��V��Rό-Yv˖E-&)J�. Hb-l�PԾ��zk���{2o�{��DKu�b�{/_�͛�g��w�sG�n�b9i���@U�'{jt�k:��e#f7t����'�
<U`i���.�<-��r6�V��<�ߞ�í�\[	�絊�$�+����6���n��Դ�I[Msc%&߶ǲ�1�ۓ\ܼ	�e�)TF�t&]Ń���W�+�^��Vo�X�s�	�3�D=lP��I�cDf��
t�R��n���U
��<��!�U���,�eV[�-Ѣy��0��h��G��ч�溪!u��~�ڽ6>Vu�QLqO,k�_��c4@
lr��:3��iq~�i��J��u:ۢG�1$�-̖�GV�-�$��[�xVHE�h�G)��w�)�@�%kk����&�� �
E���^��)�6_h�������"s�kF�7�6�H��2+@̇e�F���U]��Ryr���0T�e����@`�
�߫BF��cg�Y'��j��y�+ĝ��N��!]�8�	�C^��ur^�y������F�5#ॠ���j�5j��P�K�y�Sϡ�V�'�fB!o�3�D��<-�Z̘c͖͵1�L�f�j�����q؈	��)��N�6ІB/M/L�C e�py\+U\xL�e�u���έr��S�,�)s�*���ak��ܮ����P2״��Jޢ�̚T���������bP��9&��hb�Aݹ6�?H��{�xa����UR�Il$����s�n���$V4���>�-�����Sb�k�"���`�s]�8ߥ_k,}�鯶RV�Jm�|��"i��Y�,]o��߫+�W��Zl��ӭ��1y�iE��b��:����9��Hz���s�Z�wƓ���σ8 �R4�����55���֏�����A#���FŘ��g�>v�R�<edb�Fi����&��v�WP��[�fh�>5;I�h��8�-�R�<O?,���3�����o�t\'�j�ķ�&�2�1G#��]Z����Q0q�P�x�w�QG[��ҡ�^�#�Wcԩ�^z�%:�~�<�9�;
�Q F�ߙ�g?O�/�0�t�����6�A f�>j��^�WSɆpP�^�wO�M���'�����G/�L��<u�,&��pX
�c�34rn���sT1�l�4Ho����9Z�,��e}Ƃ`���p�������A���K�^��b�Q�F	��+<�Es��N�勗h�6c��:�K?�te�F�m]Ԩ�
����#���'��oҕS��`ʿJ�n�1]>v�x��]|��Y r<}y�N�~��JSr/NԨc*Gc���c5SR��kh��X#�����N�����9�@ϵm��\�9 ��Qøə�-�f�W����NQ[;8st��z���J5��D��u6�B�3Ǩ::�\���y�u:�?�aN,c�f�-�78�m�h�c�!����ܛ�J�O��o���=fM�ԨT�TG���Ys�ϛ�<|��5�
�Yz��Gi�M{$���^�;%!�Q`B�a�����Rl�8;6ס�<{6n�����_Km�%�U�<�b{d�
�b�Hל�^��>a/!|[�結�K(���W�R�y����Q`+N��S����ݷ�I�0�ORo:������C99����$(����D��f��6Ё�V�+�����T�w���
ՏM�c�`�V��+�h�:M�,h[����Y?:Dm�V�!ՍEۨ�o
}�����-�Li�(�#[��è�F��'�/1_� �
/���F�!N�o�>�zk��3�q�( _"��҃����G��Q
���]/�ٓ'��n��G�� �Zf5j�0Ѱ�Y�W	+481d>5�{d����4yb�6�l�����b��0�<�3�P���Գ��[�\<3HcFȁY=�š����e>Q��ǋ�i�>3{��ύ�Ƭ_-����P����
Ђ��]�h3��Uze��he��v,h��e�oQ�@W'�h�4j�֢���O�Pq�x�����*����_s���"M,N�7�H���x��-U%�H����AgJ$#d���KTik�ܹq?r�^����W܇��>�r��֌�S��Z��ʳ��5��ѷ��2G��Wɲ~4��a���W�+W�k7�������!:w�4F������)�X��l��T)Q�R�H�1ƾ;�-�,Th�\���`yc�媾�
�[,z��tN��14fF���Yl��_C�ٛ�f����e�0=M{�w/}��'�b�j+u\T�4+��ԑ5��*���G��ǹ�V�Q�P�A���~sZ�,+8ݰ�r#�����|/eѷ8^���j�G[��������冗�M-^�^:�}�U�ci�C�c����&ę�06���,L��Ï��G�|�ZG�:�Eڻu7�����<yh�d�ҷa|� -..0�����496N�����6���L�C�i�̐�>۩�P��e#  <#P��)�S�,���T��6
f�f� �BP�F���ڋ�4pb��Z�z�l6��x8�E��T�Q�e,�m��O�R@ŊO�8B��h�]̄�Y�8+Q*����8]5ц�>���:Z�r�,�r���qȍ�1ϖ�b,�ڥ���>p�]t��{��\0
����+q�/G�eσ�9�Q8��D}�9�Q�󣄆ְB���Y!�k�f`�~_֜��;�z�	9W��|΢��<4'm�vF��T6����(��Г�<N�g��3t��y��Y'������>�yV�򞨌��<ѥ���P\��hC�������s>��)�ձa���k��}���iA
0O��j��˗(_ ������������SPhp�V+���jWi�>ά&�m#�!j�V~1� O��_�V;Fk�IG�)s�/C%g�^*��B����G�[�Q�����B��� ��-�Bb��;*9����m�{��_���} �x��\��4��S�\�����%�Q�d TR͛�K1��$��`�"Z�pEq�ozM3�X�jG�ڵG׫�t���%���"i=�_���"7���^r^�u�֥֫����D��z���K��MK�������>z��k4��H����w�g>�z��Cl)���1Ai_�z������N?N����b<9/�#�Ǩ`ʪ�D��6��u�6 .��.�L6~i�Z1V��?�i���6p�q���r?;0@/��*�N^���9�����#C���郏~���}�D�B
�x����?Q�n�!��R9��(��~f"���0��zr����}�衃sG��F���5�7����\�J�֘8�E�ƃbe�I��NCKH���c��Afb�|DJ+��
�fxx
ʔS�m��B��z;ݲ�V������	Z0�r5r�ږ $�9������fq)�����8!T�6<aB],�<~���eoo@��W<3-�`E&
��#؆ۢ�Jc�W�� |�Y)���^�L^�V��ױna��jsQ;r/�u��6�W��X�,PT~��2-.�9�"���޷ٜO]ƳD˗|N��"�^�B3�#?��b7�9�g<<�1�H\�ap�Q���!��ϵF��(��UlG�ZV/����^^��p	��>XR�yKo��R+}5v��6i�����������O��*���a��WsO��u]R��X$���l<�~8��I��I����n:3p�C?�.q�&�׀۳s/U��5t`�z��J��e�5�~xչy��ģ��&�u�����WV&>�����I�ۿ�-f�/p/��;+C����k4Q���OpH��P�9�C<H���)��-O�|o�Rm�������W�Ø���.�Y*��C%��jwP�S�����n��̚>5eBi�&��Z=-���3�;�Q�+��?����J"�����&��'�N"J��ơyP	,�����1:��kt~`��^O���ʼ�B��|>��:�F�+��y�P]wl\�q9�Y��[vPD��<��-�?�/]���ۆ���b�-�p5{�� ��#��|��i07��g����J�!���z��(>s���-΍R{Ƽ2�(qU��`?)������=+�LnO���<>a�"����ή`����t�19E�Y�C{n����x`#[7^m��F&�,�����x=�E�^8�>�.˃96�?�j%E��F!e�T(�q���[j,)�Vz藋1��;����!]�k��znk��aop�	e,l�!y��ˋT1������7����������'����Ƴy��֓��P��0�O��2���"cj��+�4	�qmm�o�#6�r�T+�]�����}��(�!�!PpET
�}�E�y�ad�ShV���1fʁ������'FZ��Κu�������}��L���c�41�EtBRg�]�8���=���CW�����0*�NA�X@�� ��>{��=���`���~�<;�׽a<�JM9�FE��L�����5���;�'�5r¥Ф�rll���91���(͊���^aCȞ�dB��5����7����e����'�l�W�-"�b�%sh^�P�ո����C[����+�p�~ �����<|�>�OО�����D���^o��"�Jx߼x^n峞���
�Ėʭ�_đ��[�(ު�Zz�-VK��~�n�P��������i�ep�m���?�y��?�S�,<o<�B���bvv�J�t�֭M{G��bJk�_�d;�bM1ci��^M�7?�a��rr�c������:0
*h���w~<QlAAj�x�eB��}�Tof ���(�nE(����\Gg>B0n�(����q,m�-��>��#����X�i�N�7�i4FD�_xͨ��jz�(TŃn�l{�*%k�zE`�7�ֹ��P-�+=�l��H�����J�I��
CmW�/�C���0��D��)dE*Q>��͟�|[�.a�7�~�M_��!ao���\������4"C%lqO3�����/��=�����տ�������Z��|�@ n�ui�҃Ͼ�X-Q��љ�}�02�wc�*���x����
�[�M��o���Ҳ��43X�ˁ@�؞Z��;����C��/���M�����!tF��Sx v����}�5�}E�*1����W�֝�\���r#<��ƕ��GSĆ��a���-��ӫI��l"̴\\xXhw���5)������T1���M®7�Yd���Kϛl�"�I��Wy��|���Bf&���zK�ˬ��6��J��u|*�)�j�9��r�L��+߰�@5��Cr& �#���g�Q�u��:�(!�)��,�q=E+Ɛ����(����ʌ�Qër�\�R޼W0�"����G��Б��z�J�w�F�L���B�@�^qΝF�m�9Ӹ�ty��G�"���\#�XF�UDI� �"�sJԦQ���)*?0*Ѹ�X��&u}��*��{JP�p���XY����o;p����;o�M�bH�<@��{����^�W_y�n3^��?L��?|������מB�w(.�8������Vؤa�KNNPQ@h+Q�ɩ)�3��G+w쟻���4e>g�0�ݯ���sF���=���0B�&B��%C�����Ҷm�"���*���1��uA�_W�,�B[�5B��v�kt�s�)�۱��K0�eǎ|n8�y�|''�3`�	�1���B�idd�(�$D�������7�"�'��
����5�,�W��e|[�'l� >��-�R�ʐ�%�6�?`�ȶ��\��x ���s�yִ����G�ko�^��M��}f����~[��k��H ^?���2�C��x�96�]4��N��z\/��.�	4��]�I�7��Z:J̽�R>'��-[V��Vyg�0=����Qyx�����\��)n����2������� ���/��x2���@��.%1IՓU�����q���WYq\�t���o��ày�4B9�h��� ��ݴ�v��)��jy@_~�Es��:b�|0��@��11�'�x�?C���yj��>}Z�`K.[�V*Xp�������9������E:x�!��;:��W�@33Ӝ�B�#<�88��A��"���bh�c�?�(�i�v_��Whr|"<�S �����k�O[����>@��/��A�ڽu�-z��&�mko���B��{.V����1�~�����K܂Zk�k��!g��6t���:F��7�T�=�m#��9�zç<  ��Y4�d���CH��Ш_^RI"�G�˵�6Q�h��ͷ�ʞxoo���'	��6�r�B��|Cj:�P�������-'Z7�S�G?m��E�첒�R&7�._?�!�O�m�.���؜J�����n
?���?yc�!�P���С׌�n��xx@�Js�����俘�(U(���	~��e�� a�r;y��Ν;�#y��r��}PC:?xN�2�K[�CaB�B�^�x�^|�E�:�a|/������=��#�Μ}�J��493�O�3
�:(4˔Y�j%���XKs��fffx�<�������ڍ�߹s�6���RI�4��J4_��J���
����8!�9J���Z�<��4A�F����<J�����i���)�3��"v���
Ym�D�ZJf� �� #�;�A�Ruq�6��G�>�Q���������Ϳ��q�F�������褎��]�~�K����G?���׿�$؍�ݫ8��{A��q<s :�i���J�n�ē��*�V[7=�I�C���O�J�ֽ���`W_;���k�XA�R��(6l��y&�lbaɍ��y����hR`��2���+!x(b&ɗ��ƃ�ڕ����x�!;�IM��B�K�:r�9L0q۶��k�n�A��@��������d��#�#�i�/j��@�SDm�uF�^d�|��y�-��?�}���鞻w��}���逞�����ٙo�9"�Z��wT��!�Ç���(��$�1m�����he!S����F�����Z���N�:E���o�Vs]`\�pі;x�ﲠ5�z~~Ѭg�2��YEy#��*0!�%����&h������ɳ��6� ϖ1�s}$�y,��0Ć�~z�Ï��=�8T~��Ec��h����������1fgf�~�����n��/�2z�N�y��b氢�<kC� ĭϰ5~�7�lƮ��*&��݃Z��r%S9����H)Iv5J#=�5��b/u���3X7`�ܰ�m����ߦ���<��mO?�����TY����;t����R����K��)y�p�"���<�O<��x"�F���tH�glr8$FX�ZPlx��I�����C!�_rVAI�����K4-���2���S��|>o��l�s7�����aAp��Uޞ���p'�'����˻�C�P�V��������7^Y�+�HW���Ns���*�s�y����o����t�+���Q:~�xڴi��`}C��S2��K{/��Q4t-#�<�к)���C�4>6�焵R�UQ�|Mm"���h����۠�����?���͍?e�5?˭hB�V$k<�lP��I��г�TdÏ��7,혺-1$>y8i+�2&��Q��o��6m�H���矧�1v���psq�=��#��F�A���w�}��K�}~�a��(	{|F��F��cG9�(�+�j��~�wA��a�%�(�痾��`[W��3g���r��I���/�i�+��刮����wy�f�U��w�y��>
r.���C�
^�?�y�����Y�4-ޘ��������x�?��ve��c�3�����������_!w&9����* |mǎ�<���eC00inЈ�����(�"|��&rm:P�6�cץh����A����wJ�(̨�/><L,!�F@v�g̵ '`������v$�}�XP\�Fi�;^Cq� �@X!: %�P)2#�Z=�a�U�y�{�恉��s�tȤ�l��d06&&����."c���ږL87܇<��dL 'B�H	�!�54���o�(����j��6Y��K�sf۸�0���e##����%���
��=Q,��ᇲ��{�p8xdd��?��?z����y�n����g�g8<Ξ����û�K�w�f���U����qq߼��|߰!���cף�>J{�`?E�ܺ����.�$%�iqɣo�˞P��	�V,�k�g2Zwu�i53^Wr7z0ُ�q�:���aBQ=|<m��~�F�w�vH�
ڮ.֚/��o�B�VG�2��␌;4>��(��������C������u�\
,Ա�1��0xu8�֬�3�;6p��tq8�@�Fp��"4�漡 ������6TSߠ�"���Vi�@ IC�s|�8d��p&�T�5�k��7c��l��"�
Q�4�v)�nU�����dT�9�b�ȹM�۷��sꉋ��7R�p/(t�����d�4>�H��4!H����w�aІ�pAL#�r��v�UmլE:�rj�c6�{�3�|8/M���\��
3�T��/c0�'�����;n*�[h�p�5s�hz�ރ�g�.:}�43p�H��ݻhrbR����+�����k��n�*?�nM�FB`���l����Gh��m�o,��-�G��������ݫ���(�Uy`7ZɅ˼����_��5aHx݆�^C�`f;X�iȐA���GM:ySs��9 E�8L]m/~B�RA�����9� t��ব��:�|y��K�͛7������K?W�\��i���,,�h�R7�7��o�` L�,��{�N�<��Ixiz���6��,��V�
T���e�V�\��:�<���(��K���X A1b�P`
+o���}�wzz�:�o0�(�D�Q|������h��g��֩���r˖�l�@���^�pY�k3�ŵb�y�����;^~���C����'$
���[W ���^X�f)��d�����V\\�����r�6B�p�[C[nP	��R�x��o5/�F�\3�eb�z6n�Ϝ9M]m\��a��#��[�;mٺ��#fc?"#�葇���{f_AH1t´�{#������sm^J�D[\)�!z��/�\��XZ�-���FKz]ż��^#�G%�&�[����`|��B���$Qw`�v�x[��¸�1�ܼ�����h��}��Z^\d �"��g ��gjY ?�&�Q�%P[���bphh�K�i���4��ܰ=�����4
���K̢��� �\Sc汰�H�����S�~�o@�I�f��p���t�� :OQ�^��r�Ê�쩍*Y4��5Fĸ�8D��G�6��,#�<_.�u���>��{/��o�&��2��?��l��K��M�u�+�1@2�y�0����/�
�y��%|�{ߥ���o��FNh��@��;y��M�榢9�,��z�N��X�w�	pE��1��_5��F1��Bk0t�<I;��aX�&J�4[�!&7BگF(ޝ�����}ū���'��e�_��?���z��W��8�<{��z�ѳ0�f����~��'>�������磂i��jD��щ��=����;���/��/=��V�-���V�k���|�җ�{�m}ܘ��YjJ$����{��m��F�}}XYM����6�8d��"�.�x<�it�i4�l����B�(� ("r��pվ ���CC��S��#�����ؿ�È�O�d�X�EQ��7�
�(��,��������0
KA�����SO?m��\4��_}�U�O�D�/R{W�6z򳟥��}�쑋�X.1QmGwU��x���z�����n^���i��������äو�E��� �0O�p��zg�0s��^�p��hP��  S]IDAT��(5�l�ss�t�,<0����Ƶر}m�돾�o��t2s��F=�Ì���6q��ҁ4&��aшF�5��[2 +@ԿJas�g&�=[�G>p'ݴk��Й��tedn7�����h��-�ꥁWipx�jF�Ȧq�����u,񲲞(%�U�q~�k_����7�G�к(�7^��h���_l�.�C�(� ��U��m��(�s_r�1]T���� ���"��[o�`oʯ�ƪ؊sYn����b ��{]b�dzj��t��-@�a�(�'Gd�J�FЁ:q�ǉPa����m��`������5�����
|����F�3��$�U0@p�J5f�i\/	�!W%
l�'<5��s�( a H|{G{U,:˭��Wt��w�����s���6�O���K�o(2��	�)'Ze���tӞ�t�� U�*7)h�}���G�?��_;` 9�I�d�@~(��0O��Ν;ǡ'4�	�tn+�e�si����ꁸX��B�͋�	 �ŋ�X�B��Я;�z}�; ��{������B��5{_�Na�7��h/��&��=G�߾��nl�o�eʇ�+F�թ��H�ys�M�b=O[�z�6u���ƨ�s۔ڟX�S�o|����ZC����;����M.N�D�	{��aU^ú�_]�F
�7��Ύ.6D���䅅�/�~
�&/-1nt�m	Ci��w}�8\o�I�V�X�;Q!�hª-���
$$��b�Ꮅ��v��lڴYpC��p���!�	i|�Ĳ�/҇s���;���_��y�rY�Q4��B 7�e�)�Է��=,�	Y)�+Q��(Dl�r�_ö��b显G��|���P�{��G��s���9Hl;�:��Y<�3�'�le�
�%����x+u��pP`��LcEd��K���[@�5V�>;7|�����^+\[����7�w��?������IƂ�Q�و���o�c����ݶgݴ��() 8*�˜C3�F����j ϟ8A��;i�;(��E��&iѓ�13Hs�Fs�^�[X�����F������EqC��@��'0V8j�얣�Ѿݼ���'�
V�}����|������)6ُ�������ٳ�-\�}� �p��z��� ER{����|�2X$�4���k���M\+"J��~�K��^��U\xP�-rW8w$Ng�C�}�-�p#塨?�q�=�!�S��u�\��"2E��Z��F��ic���{�P�
�����:�n�K$dF#��q��dm�Y?���Ee��L�W���'/&���_�x���j$��.(1�sK0<�p��L��د"�-
�*6�"�J��#'J�-��ِz�2�)S[4|�����
���0�F��ˆ�v���}�0�D��Nj�4��SE�f��fWz�-���"��q�V�����{M������br�0��Ӯak��������2;���-9�;#Dୁ��G�]�v��jS��n�XbgM
l�]͆�Z?n2���{0�e�5d�n��M�����{w�
F!�9��#�etB>s�,]����r�婥\{t��X�
;�p@������jQh�p�x1cD��GA���N'���8Ma1�bcԛ tjA�ϥ�!�nx�����Qԉ`�Q!T��R6η����#VRZ��ِ�G�H��3nc�P�r�������d/1��<ao)�)�� ��:(a�GG�ޞ�(�a14��24o΅�����B�z�M�^�t�C>���+��Тg�Гa�"E��P���m_o/s8�5�uv�a\�u�9�JU��˨�����]Y�;��٦��s��}�!�e�:e���87��;*g��E�4]Z�:���u��RdOnn�DY��|G�*M-��Lm�h3�ZA�%�C��*)�GC�<&U.Y.��\+�	�@�Q����`�U O�{ ���"0)0��� j*	���̳400@�NО={Vui�ki��{�Շw���3ֺʾ��(mݲ��7�S�`�5�#�Cp'�t�� |�=9rdi輛[QT���^�؏_�s�)8$���ķ�/:�v&U`�����[#�X�@�!�w��I�\+e���SO1�[I���j�&��~�Xh>���p�Q(���"� �@/u��Ebqi{*q���Nc�gPGg;q^|�;�f���({[٬/�\3����n9 �+L"^BaM�Yo��v���֑���\ڠe�(L->�b(���3�{���@T���@�B��~c�΢��Gc�2�7T��
9�cEUk�p+���1��w�
]���F�Tz%�܌�e>*���8�ƌ�W(�Uhe���$�-��Ú������`�1L�y��מ�bN����TQ��cšx�g��l��g���ĳ��Pw��(�S^�5gs��`��BYKTA�r�B&o�\d\�|�]�F��1EW���	R�vxj��E�j ū�tc��7�u����>V1\|� X�D��A��<,Pd�֐�<�J������T�	w�����c:P}���q �si_��/ҷ��-�h����~�����������J/%!���>BtPr��̞�5�����$Ǳ��H�//��
�/鍊n"%�%�}�;�!]1��3
� >k�Vg$^2,����K>� }�_`Os�pA�t��z�k�� ���R��[F��n��&���>o~�Lcc����1ÿ+�|�	B�����P�B}v�q��SkHZP�\@o����czf�f�Ok��9�u[75
\���qa�r��Y�(����/:5+�w�F"�B��})��I��������WH�ku����Y�칳4;�1[B�ڕ��-lg��>����	�A��"N�\�~�=Bj(KU2
���5+��=�x���!z��[��n8͗��T~A�C��~����K/5[h�p#�q!�4���"s_��UB�+��؇$���}���("��K� ��)���k�IDJ�DN�̋g�����g��PcE��aǀ����ыf��i:�y>x�M3k���SBZ�퀵A[¸K�?!�0(k�µqU�Ѝ��h��z����>��$�]�#F�]�2�����s�������`X�,�G�LZ�I6��~��bܢg�8^�|��E�"�����<5�3��p�k�ȃ!�/H?1��2����B��Fӳ?q�8Tx�1`�6o�c��s?�}�Q��׿���/}���-�&^|�ǂ���a�뗾�kl<~�;ߡ�����M�+��a�<��\OH�%yv��V~F��a��U���4��^�,W'��[�4����[��ĂGv�T�Z�||�\
�*K���p=3�g�Sy���n yA=�ś��h+�N�]�z�K���<@%"� d`�Y��9���kSԢzu6F���J��@Xu=(Gq�V4�3B
X=Q�
[amk=T��"j�Zx\����T��~4�ﬨ�����.a����M���B1dpjn�5$���[o��'Or��ǵ_�_��1l'e�D
�Yn��eғ��P�c�'eg�8�y�U�C�k�\�o�Ia����)�#�|6m<-P�e�u͚�����T0J��x_�L�U�)�-��Qe�|٫��	����~ݾc�7�0GO=�4}�}�y�R(�}������ɟ�3�<���5ƽ�!v!6�$w�p8A�U�%t�3�_ٶ-�P��i�q"�'��kW`KXg���x�rÖ����H+����r:�jh@���WƉV
�)�
��p^-���2Cх�)�E���#
+ǂ�A�!)��,z�`�h0��<���0�^f�0&���a�e��v`���\�Gv�:! �l�0S�\�V�.��!,�saD4��i��J������y���`_`QA�3�b �&���1����ʥ:�����YPI6Z%�%Z�M��M�D&_�
±S�
��;�7�`�8�B!}EJL�=�߇�P�YVn��*���߾�6+Fy!�/����]�:����c�t��t뾛���G��Y:52E�Ǉ���4	~wp�=J2�����uup'�[7��-F)Η��u�6��P��l2�B#�� �B�05N4�\W�R7$�3�G��g���7�E>5��zh���Z�ʫW`���_��r��I>!4!`���=Mc�'�݆�{�����2��4t��r���Re�]����3y,.�G�&�TP`8g�؃� C8���L5�e�߆�M<u��%�=^���XE��@�XA�ª��N�:ůK�%%	~�A����`��^�BhG�9=�-�aPz%%V�R@&fM$Ĝ�G���J'��.Y��IF��zfPR�P
�<�Kp`���)bEm�����6�X�ֈ�Ii)�z�1��K'�:1�L��7C����襶n��(�Y�"����6utȊA322J�/�b�f��u���@f�+���u#�O���ct��9{��y�L�a�	�<.�ڴ�0)��mۤ͊���=/� �̘g��9�=Y�X�I�>+	���Ts}
�=���+0o���۫�u����p-6�=qhݗK�����@!���n����M�}���7�
��iQ)��pC�~��c�X;|x����ٟE�T�e��������M��g�2�H��!C\(�bo�9},��y�0���+tl_*�����!���cT[(S>+��n�;�@�5,%�S 	C�5nغ9 Y�$5�v#��&��<�Ud^���u�%&5y/�sK��(�ii��f��ב�\�Tܓ+OA�)��gl{P��b���O�%o�ں�H��m�\��bp�R�<��166M]�N��L�����-��2`&G��u�J`�y�s`��W��������K��K�hl|T���������i�/�(��l�\F�/6� �/�������9�������ԯ~�WIk)�sW!/a	[�����k_K?���u���5ܼ�*���H7��� �@FK ����̙3t��1� �u���*�2qQ��[PL�]�'��<��o>>S~CU�P���G���0�| �>-�غ4����a�Y�u�>�4�Ŗ_�q��Ǐq�S{[� &r>��@���((�;�����9C�Cy��ą��ә���={��o��?�s������ǿ�}�Mdš	}R ��s�R�É�ۋ�SJ�0��61�A���ﺛv���
�����λ�RDF�X�������li���*-O�1߾'`�:	����t�.T6�i�ƼԔ�x�ϫ����o�6���>�����,��B���(��_z!#9�Z=y�$�8���v=t�� ����W^�'���;A��C�hM�;�M��+����_��^{-�*���w���ХKf�F�o��CNmC��N�1����o��:��������n�G!����ߥ��u���n����W^y�(*e��2Q=���-�OxJ׫�8n��q<͓��9�<� nb�%B���P�$x��9Z;��Y�T����bgrr�-fP�@�A���gY��9����z��H�@��t����f)�s_$=?rX�_a!����-HZQ�KZB�ɧ�6�.<��|�3|�F�^eb�E�l�!h�^�k��B�
`S��J�t�X�����f��
���?�aڿ�V>_t�������pVB��.zN�+|V�s��I�B�v�g�C�����86GՆ1x�ݔ͘�o\�E��������졛&�Wgh9G���eYjڑ,t}Ĉ����GF��>Km�܍!�I]�_x���.�V>�rx`�iVZzaHA�Ã�1T��#�!��u��l玝��U���ӑ�rÅ�c^q@�yq�פ�n��r��*�p�����s���E��`�Cy!w��N����Hr0�&��z������
�׺!�
�\�������yCaiO-�<m��PFz�EUj�9��e�Ŷ(�EN���C<w��qH�5"f�]�o۶��I�'UQ38Ģ<��ؼy+{jX��CD�g,1qJ��_�N����s�0w0s�0?�4��6�g��v���ؒs��C�����p�s/�c�[K�sa.c��M���������ڊ��"�N���\�v o���²�5�)J̏�$���Ȣ�%��f����B�A�Ec�亨��)[졁�]����Ԣ�+:�v0�>^Õ=0fZ�/5h��
�9wV�|C;G����e6�Vb��(�G=#�׻P�1��W)��GLx��!;����Fa��|yi`V����8IM-�KE��<��X�P�^��*&�*`5�Pݴ�ށcb���'"᭞�6�<z�(+�V������*�t(�i��s����a!/q<xX�T0sr�z�k�|�]��Ҳ׻U��ň��#Eesln۶���U������ѱ�U��X�V8t�(xe��h�i�Pq=7o�le�=9;�5_����K8�J���0Y����VhI٧�ӧ�hP����8	x�σ'�����8�	Z��B�΅�t:A��/R�^����Q$@$���()�w��1�s�lX3�-��\t����x5!��ZoH�4��M+XH���e����7��[dk�m��x���?�ڽC�U������Rq�'�WT`���*��5�����ڇ�2[y��PL��
+��F0p���bڻwo�w��n��T�!��CA(8��n��X�e����r�Y��ض0���A�����%
��0���Y����;:?x>��X�H�C(�����*�W�`�U=;�}�vӧ>�iz������
�瞧o~�<GU��ǆ����*�p�p�#������L��_��Sd��iR|��B���|?VXAB ���ja�[#@�����=�i��A�B���#,l��7ه��q�*Ȃ5t'�ReH�š�\+�L����̬Qkx�Pk�"�A3�
�Aܬ�����
!D��*��[^��(
x
�-��͐؛��c��og�_�ϥd�1~l.�1�Z��f�׷ =|:I��y%fu}#�����î|��Ʊ����;v�`��-vl���P�9 \�0 &Q�*d9U�ڲD�NG�q���e���q�=�BF�L��ƛor�
�pl���O~���}(QS&��ϔ;��@�ݵ������λ�ΎN�	�\3��!<](1QJz衇9A��JUH��z�����¸^
�@u��8N=��g�F~��9��{MI�^�������5�-�<��ii=�\'��/2V:D�sA��G���W�T�PZ0 �����F/*��Ht�����8O�Wrg�P���,�[���
%~s�,T�MT�7��(��E���OY��@���$O��J�~�z3^���J������-{�k�HA��<���F�S�lQ
&��g��k�̠�aq~N���*/�%�i%)~}R~Evc����y�J������h��l7:t�B��i5�
��q�
�����m�6�g?�cen2z$Ö�/��F�^���_�k:�<'��rŤ(D�	�E�&B3�;t[��:��?���O�́iO1m�	�`X�𬴖
!E�l^��v��0$�����7+i4�rCN�51 +�?.P�y(�%+ߥ�8�E��n��bD�ZX� �Å�fV�6��K+��X~��I�A\��Lm�����F�}�(t���10����6��E��Iy���`a���O��4B�(�φ�B��
�)���W��t�"aëJ\��g��p4���q�Ǒ��|@:5���0n��+���Ac�4��a�[g3�)��*����vE���jv���և;�P!�a1rh10�p���V`�S2��+RB\7D�*�H SR�i�HR���y��4���|@��"N:}�4��TFF \��ECai_o�(�O���;ȹA�p��B����J�5=��l�_�΀@�g�;�����߿������eL�54����	���^>~��g��o;�1�xq�(.���n��1_�Iu����F�^X[(Y=0��n��x�r����w�����s\s&�YA!t�R�l����]��f�5��J'���` 5BQR�Ƅa�,5 �LA]*���Ҟ#����桽�t��,�^"Bf��-�����8��k������a����䉿%"�I0�03��nZ��>��n C��?>�Pd�D���[�p�r[�e1�>��n�.k�����!Bx
�ᆗ�o� <1X�
�w��ܹ�h�DcE�V��hH�˄�#�z�UY+PE�Ŝ�33��/!4 ����>��G^�em{{���3gN�B���[/��\���t/�Blw���Ea3��Re���RWg+��i*
�:�����GO<���PWv��1D�EؔZS���qB{C�Sk�z.��ja�*P�s뭷У�>��<` N����d�;�2��� 9�0�5��������|�gÈ��E�P�C����a[�4�)�w���r�qK���{=��O��n��L�N;I��{ﻗ��_�U����?�:0�C^ͣM�7�5���ƮuGG��x^��=��4 �}��G�N,}*kV`�B�{h�
�鉭���uPh�T��e��ӟ�4�Q�t��\�p�_�@�iD7���I4���ϦH��� y07�S�q�!7�`�o��6��6o����c�ya�BT+��aÌ|�[���QxQ�����B��@~�YչFm��y�����鮻��: V)a.!>b9r_��c�TK
iO����_�p����0�/���u�φ�{$����tA5с�w�F���\#�oo���v��2n���kٰ!d���a�M��Q�6x}B䮸�ڋ�	��"��P�o+BPz�i��X��J8>�����
��,�c�:�K7n��F�E�L_�BV��+#W�z��i�����4�СC��B���_�"�o_z�E
�aj���`CAZ�w�r�q�^ȟ�5Z�両�g�7��ֱ6L#?�D]�aBZ�2KGF��l��ו��s �����t
�޿?[���{��G��,�c)K|��#rOxp�ԕi��T`qhIl(�F���*'�,g�:����-po'<ع0C�=��6�^)�����2��sϱ���~wtt��Z�/q-�����@N���bb`4̜o�h||��.��P�T2�~�����d�3|y��?�F!v��y�X�����Ϭb��Qg�!?��Q��ste�
y��顳���(̜��J���4\��#A#�PS�!%��t��y�oC��j�JǄ1�5��bvf���ٳ���c�4[�c>��0�����;s~J3���F5�C�4n�"^� '#����y��lCRl���i��	96��$e�On�ڄus�����ߞt��r�&�&�7�ܢet�6����KL�u�S����Ҁ��ٹ{m��@�|�z��W4,�rP¡ X�s���*�(Y��ȵ�iG�FL\�fO3lu�õKx�-P��%������j��{��[?���p!~�x ~�a��Y�[M��>t"*	kE.��w%�E����2a��/��8�߆Q�D��U��e�i3��n�"��u�)�>��� <1�3�PQ��{�nn6�L$��(�e��zW۷m���4�|��%�*�ǄDX��M��@K(?xh�p�8�|�#F�M���(��-�R#�ܤ��@(7(U�XX���9I(�j��2�K_+-�p]K���%�6=��GF��>'g�ٮ���8�Z,�FB��3��C����~wgN�Q�U�<R*d	�5���2v-��LÔ�(2A}ʜa5�9�Qvh��Ϫ�<ڍ���tY:�?���t��m���<c���n�}��{z��Wh�P�70p�n5&�r�ʢT_B�%�P�6o��D�͆��t�P"��pp:T*��F�������[��Pd����F(%�u����	t����,z"u3�Jhnn���l|����I�0�0"���i��W�#7�f�d�=<2�H?X���y�/�mQ������f����Q��bU ����ix�8o0�4,xb��hX#�SaD��z�aU���|�7������m	�ڋ��b�F܁`u ��eHDM�.��<��Q$J)�ߋ�(0��VW�Q_�N��5W:��ܞ\�O�^|<��ye�(��=!0�ј!+�t2�� �����u�o�X0�I���gϞ���~���{��?@/��2�s���֘XHP��(	���s�[Ѳzh�Y��� ܰ|l�H�\�ܸ���
��m�wh�sU(���>~�c��-�f�=:�F�؋�=]4�Y�Q/��J�	�`�nD��lG�	�&�Xn1�A.X�$���CX��L� ���BT۸��`a��AQi��łg'���y�ܶV��(�B1�!�6�H�M?���d ����֭[�ST��dB\����R�����K؊�u�hD����gA���P�|�^��<��$3u̲�@q��j8��P'𢧮���j�yR*_�G:q�ZD�{4*����_<�L��c�XOƓ5φ��7�Xfinf�C�~����o�}�Nڼi��T�s����!~��t`�s���L5PZ7�Np�,����UDZ/�ϵ�kz���
��PP�}q��Q�䥷�U��>sw��������kk��j1��Ei����
Z.V%��S�Y(��QҗK��Y6���bp:�B����`�<qP�'N�`D��܈5�+���J���)���,�LF=�{o��i˖�@s���e����-[6�8>B>n(�o�� <�]�w1	�������J��+st؋�Q�Jț�1����{��wq��QF14t�!�����&�R�P"�o�����,�j�:?p�Neh}��(y���x/���}��*~�1q?@���*c�P�`<0����;����_X6���@q�A�Ҍ'�x���n����>5��;?j?��������Ç������~H���7��q.[�
�"�)t���@�P^N��������yICNKU�떺�e��po��]�[�}�8c]q����u5��XMC�1���P���[���Y�P�̄!�fc����?�A�2e|�.Dև
�V�rx�C2�Cw�$�%tc��B�E�e(ۖ�\�e�3=[�BH\�e����ill���{h��M�X��� �u���ފ�2���Adsf����;詧������p�C�%����Y=-	I��\��ށ�����8G�5 �״�X�d�J�^���xׁh-��
���ٜ�y��Kި�\O���B�k=�gߨ�<5*��7R�!~@��,��S�^�2�2u�yzT�Y{��$ˉ�_0�k���c2�(�G������*�^8v�=~������zf��A��;D��g�y��:c��>��O1��KН&3���~t�ٵ�k�ㆅ���c���zw��z����e^%���MJ��lN��xx�^dui���g!��gO >��o��ߨ}Ӽ��m�6�Y��P!ZQ�8ŵY����w�2� 6�f?p�Az��[\���5�e�s��offZ��Y�H���={x��S��B� ��.d�B���i����8�����{M�1�Sl+��Q-e���>H(��CD	��a�I��^��a�wʝȊ~U�|�g!�UE����be�✟���X�9�V��zw����h*���%����`��(0(�P�.�iD�g����H?7�5fq��o�%�6Y�����{�!_whg���r� g�']ӗ���a�� �<4���[�J���XV��S�fk�i���`�&�l�/F_Ӈsbb�n��:sf��Ѱ�+���{�3(�</��+�� ���~��M��X�Ԥ�Њ`��>���n�f�Y·��t@�Xȳ1� d�圠T�#Sa��!��)��}������}�М;!�`�%�0�gZ%��,��5���?<�K��x=$g�`֐���cc#�|!�E�)�]ڤ�0��!��'�9EB���\�����W�_q��=KE�}Ԑ��mC�QD��5�m-�M��9��N��YZ��5�V��MF�Y_܋���c�ͨ�x*������W�ǥ�
{X������É��+*���6�!���%���7�P�E�����D����}�c�P�yp�d#@��Ϳ�b[VA�
�m��F=��|���i��g����o��BB�l\���~���n��;`�� ���_d��
x%PnP�nG�Y&���^[�����z0���P`*�0��Ā��s*���[�cA�����тR�1@�Ӫ%�U��"�ƈ� ��"�0�||�X�Ԋ�,R`VI�"����x� 0�z�($���l䥥�9nX�ńpH�Ea?��p͵d���эd��;�T�XCo�Nv5�(���5�֕�/�H[�7r���+忖{_!�@�]F�A�j�.x!d���F@a�- BV&/#�>@��Tţ��
��i��}��N+W�3`F_jm�=��z�r�g�S��͛h�-�lk�s������'�n����PNh-���M��ZAO%��Ы@�c>K( ԧᵆh�ֽ���q����:��&l��̙�
�����ѡ��[ 8~�G���jpjO���
UW�f�9��� �U<RT��a�[�bx����ߢ���Q&2&�o�i/|]EF��6��^�vS�d��c�3Oڟ�~�5��S�On_���80��g����۹c�٭:�����KΆ�H�_��݈���M�D,�,�1�=�}�5�̑
�7YICՆ/�@� �hUR���C�Z�]w�4��6芋]q�����5�^U�eI���ć~�@� �da�z�L>:���P;IglAv	�G#fň=$)�������cA{@�1O��5�C��:V^aJY�߳a�P�S���r��x`��u��׌B��c���z$ �ԍwZ��]b���h��A���9s?dѴ2�l��Y��ڍ��5l�dI�P�q��Z'g�bXC!�^�2m[�A���P�tf���C�+�A��Bh;�f���vÅ��Q_�H{fꌶ:Zv]���_ܑ���� I�;����ܔ�s�^#/���B���5���m,̶�I� ����g��A��X�6�ɵnA�{b�C=1>��OjӦ��Bk�W�ݚ�v�����z|����0-��2�Ж������V+n�9�k�Zc98��v;��p\��8uZB�6����� -����XwR)sܢ���A�ބ�uX��sQ�Z���%cK��ge���Ή��ъ͛635TGW'	9�7��F����oa�gP=�����6���ѣ�&��P^�_W��p޸���r��U��wV偭+���y���![ P���
�iA��V�hy��<�$L
��О /�;�����C�	y(� �<(�����#M&E+B��;���a�
���+��<Z��'�+!�T@��"B	{���x�����ů���'�*����C"E�R$�����鸌tYV!)aJ�γ��)��婔�&=�T8ב���s�{�������W^y�.^�_R8J�l�S�:����y��;��P�J�2oY�x��e��
F�eP�t��P�cz�e����@���;#Oj��{2�9tv��w�N�>�8u�d�3s�t��&#~�ɏ�]w�!������Ҿ�n�<�D�n�R�jX�j��Nγ��;�H��uw��������0`��.�cW����T�\�xo���>���Z՚a�5i>��)���+�DA��$��%��J��9L���QB����Z��(��K�A�Ӂ�S����(.�������T�A0���ܹ�FX�gE�s��Uz�'?�N������y���ۥ{2�B�x P�����g��E��`o�o��!�R�xn
 ��¥�"�s�%�B��ߡ*-!��Z|��j�]8/j-s *����a�!E܇���)�*��P`�\>OZ O
�W����f��:�	��h;-v��BWo�p���mn1�'<cl��8�H^Lu�Z��c{�\f��s�ŗ^��N�}�!����[��Tj)�[=?���Br_܋�^ەj/����/�@���N�:֔�Za���Jb��}����+���j�
j�ʁ���0&@� ��x�!\�����׿�W��<=�@�Έ6�omٲ�(�n%� �xq������?�!�� �����$�xv��'��~��1c=�8~�~��`<�<<�©{��^z�ez���Xh�%��x{�	ñP
�$��|�6|���o�����~���?<�����u`|R�-]�#�vCHq��[;.���YpEݢ�t}cd"��{����|��kF���ѽ�⋼��)<g���P<F!Hg��uFB����y�%��}9[?�%:�b�::l�k����M��5��{$k���t�(�?<`��<���kܶe�����{���V7�]z'Q�ɺ*���QNݽ�t�����q�Q�����ǎ��R �Z��%��u*Z����t���+�h��S"_70���U/�e�I<�^�9�v7+�x�_;��}nW��V%!�k�����hK���-�DHa8��r��S��3
�d�Ŗ-�}C�۠��~p ���po(�j�̔O��/D�B�x��;�x>�$3l�l�7�o�;g��s81Mڪ!#���[��$���� �|�2��捘=�͍	�$��<��"�H�I���������5<��C9��;�yh�a��g,�;�wf �;m���%����*���x���$�ć._��M�!G�)���N{v��ck뙱�Q:�V9ccQ��g�޽\G��[T~��U:u��V����%����~�s`�A��S��ܱ}o�{ �q��ۂ��q�`�p� i4yʘ�0�@A��� "�84�o$,NF�@�%�i��U`����:������w��"�Ta`hx�_4ħ
����X��I���\�}h�a�WHr������A�lV��|�A��������U�!W�f�����Ѧ͛ٓ�~[Iԝ����� �^�%�C�|d=z��l�(�j�ɂ����!e�%i�7ev�zͩ+�,@%VJ�K�u�۴��
�eߋ�eF��r�Y�eXh#��e�Ȣ��k��9P��cZ){t�n#�u�]L�0m�(�B[�&g�8D	h;_xmw�y'}�7B���SVw5�Ope�}Ev�ۻ�H�_B���Fn������c�m}�_���?�[���{�ᵘ�������Ek�4�@��PP@y���z����z����N R)�*[v[v�D��P
��m��֝����0�F0wA� ,2x��9 �Vv���L��Ɗ.�h�T'�U�����p�o~~�[V��Gh�FCJ~�R{��yx7��)�Ռ�P>cC�hP(�h��<�߁B�%�HpJK{y(0�'i�?n�^��$�c��< � ��Ä`P�ݎ!G����J��g��R�V�XV��K�_`�QA(z�'f�Q����
����s"!XtԾ�Q�x�P`��`��*����\�uA^�K��ɥ�}�k��b���yj�ׄ�!:;�6�'��҆66�b�yV��K�T ����{i�QH�:Sc�`�������x�C�o~��z�����O8��ܳ��������U�:2s�xFЊ%&���"n#�M�D���k�L\�*��J��C�Q���|��X͆��o�G��Os 
(_X�x,�Cz�f��O�37LD
<('O�d��Q\/��#���?N�O�BJ �ݸ���#�x�~�����PpB���*w�!X�(im�z�* U�@�6,T<���o��НZ�؇]�~I�Q���;"��x �e��A��Q�u[ ��E�6���S�BI�VJ�����V}b�� t���������5���Yqq�. �����Ф�P̷^={|���<aC9A�*����ݏ�ge�X�8'S�8�_���1G��o�N����g���|��7FR�����nΟ?G���oF� ��Qņ���r��H�yd��q���?��ݹ��Ք۲��8?�G��-+�43����y�-�@��XW^����`�f}���q!�(0�g?�Y<�>��Oӝw���B��a-?v����N{����u�{�9��y���1�喛���Á映���׾�#��nsl�4��z%Ou��<��ssJ�!�IJF���u?
�`�����sQ�k+�d��`�}�R1	:�#יH�6�}x�+���;��s��?o1���Q+ Q|�܁X��c�ǀ��\���e.�c�Mcsk|B�\$ 
�|s,���{Q�MSA�%��m�������c��0�^h��z���xZ�������h�E��%�y�֟�t]s%�t�"MON�!��F���]�W�ȷ@#�С��ˆ�e��`s���������P��>X��C���k��Q[����&ꦛ�ѩS'Y�l۶��?xo	OV���l�D�@	xxh����I�\kVY���z[7jh�K�	�9N�;
L!��y��Z��_/�7o��n��)�Yr��L;�K�" �y\;��Z�T`�xa�E��u��5K�=aÐ��
i��*�G�/+!�ZB������i#�ӕ���	�%?9�q3�U6P�=���+FcL͗�T|� l&)N���0�A�����9�T0@y�ڵ�s]h8	�r����i�F3�QT`1���� Pb�|����%������	$�|�+��ױ�2Px��A�	��VC�Z`��ʆ�-�U�'a��sn%X[�����sX��z=~+�I�<3�V�P0���\�Yԝ)��B|������p�G���������nF�Y�_�1`�f�?���y����;�)�,�G��L�L�ҫY��APąӾ7�p%��V\�{w�EĭH��J�FQ� E\��f1����GN�n�_�ɨ�ʬ�����iVFFܸ�Fz�{��ιS�e�����L��8)TB��?�-!��R{�ߢ�V����P�@���~�ސ��'@CAQ]`���ŅR����իW%�f�9���?��J��jF�$� �8q�ګ
��nP���ѕ�s̈́���XQ�����d�Ѡ�.%�X��P�XM�W	�|�>��rq���wu�Vu�L^N����X��5��2������z�j��PP�&S_����ϟ?O��B�KL'18s���M0�*�g��n1G�>W�F3,4�����Dw�BEWp'�<��6���W]�;t4:��gk c��kgЉ�'��������f*6`uP~��ʕ+����/^��\{(
�B���7nTʄ*(%�"	e�Ju�ܹ��ѣ��ӧ�&���)����iś���~ɫ���4��n�9QX�^J2A���lB���,i�G��P'ʙ��"R� q 8iQȞ�Ms�$jHT����}��o�!h���-	ـ1KL���e:�ͤp������4܇��+�[�}�;�����&W��t	P�Wd!�!�Bn��\�SjE��q=�5s���A���:���.��&����z�,B
*��d����T���ZY�b<e��u���tL�;��>[����������+�
�q�c�J�ٔ�A!\ge���Ν;	 ��+!,�~�!��J6�k� ��v軄(���@BA��.�^���X�_�z��e/'�3��e�u�; �0&���+�{,K����6��5�=Jmnܸ1W��V`dsNI_`�u���=�*��eZ������x��)��D�FU�![�fMR� =����֛c�ϫW��r������\��2'��|�8f���U�Vf��O��qv_�&/�d"�M'ҹeN u���i��Ng؅��lD[u^i���2�n�j�"� Zg��\i�Nb5n0^��H�U��BBh�8GU�)K��q߽{����j]N �֒+{	� �����>��@¼�=��u�>�ۥp��x��<��J�0�E͸��� ?�m����1��9n���1N�բr�"����]Y�)�$!U��f�d2�g���II�&$�E_ ~��3�"�x^�6?��Y�`����y~9ݺu�z1��9Ɗ��>�XH�R	�"�6��2�����jMa��Ss�8���c���Z`�,[�%pt!�c1��հV�߹�+�l����+R�X���ݻ�}����Bt�2�?��_�N�A �"��6�FL��͛���1 %��E���ٓ�ۊqA0�r�b�z5@ ���t�aq�^E[m"Ƶ >;w�,8�@Ǵ�{��mR���J�� -�q���Ey�֭��l <�����W�U��y���0���d}��g�߸%��3@^�|Y����i��E�Xo��cQ���%������XT�b��7���C�q�'� 6v��`u�mS��a��\%� b������Ⱦ|���c<Ķt��D0��ߓ�C��{���+�
�q.������H!&��D�CP�Ϟ=K f�-Kڡ|�Elů�	��l�b<�~r�͛7'���p�	8|� #�1�'���1j}8��I;����`˖-i��L� �� \~l�Y�qv+�CU�h�M�Ыu(�2N���\HX���1V��%i�>�E[���V�si��\s�b^�c5��L�/�����^}���eZ��[q�z�r�d��'x�6"�ug8��V�C��a[����^h6ZZ��N���:q��~�m��s�.ȀV�@��tK�7�a�:>��L�s�F���(,/@E��w(U�+�/W�֏D	c�Qg��$�J�:����qO��(���i[r�1.�խ[�V��B���K��&� !�0�%9tGP,e=�n�D�9��$�K0�9v�t�s|&~�o�v꿉�_�~���c��� K�O�}J��Y����۬� �놖�%cmh�%�f!����!3YG�}�2캦�#���+�X��PX���[h7׊��3������M�QD��p�b�(3K���ï���W��(*�70$.fQ�I@� t���EW��3����u'�6���t:}FGN�X=e1e(�5�H�>�,�ZiY��ɨ.	"��f�@:J��"�Zѭj�sdZ������'ݛZ{n�!St�q&�qk���d���S�8����UK�De��K�Q��ժe�y��lD��h�/&���EV�:E=4��2<尕VF�&%�C����)n��҂�
)�R��u����[Fu7U]a�&nD��l�Y\�����Q�ڙ�2���,L<ۗ�7]��a�S�͈�?��,�t}�e�_�
>&�Z�q���c>`XbT�99���1y�Z�UJ2�lX�K��f����K�F��2����hey�� �<�XU:�*1fم(@Yk(8�N�L�p ʖ8��m�1�Y4�U� P�D�'iD��B�ⶴRd[rL���k�H ���Xa�1�h�r�yq�:8oc�L[�L�y_]��4>�-��Y��EG��*�F�.]���;��x�0�%ֱ����`��x�}nQS0t�C��v���]�ѿ6Do��/%��d�����b���V�@ѩ8i�ztT�WѢ`��U= au	XQ�=x� c�Σ�Q��̙3��V�҅���8���G�%w�F)c����\!�)��V�М),���vF��t� O�,@��冑�7�-ON����ə@��]�T3I ���ݛ\��t
�(o��$i��^�<��{�!�*��g��|Ę�&}�恵��2��1�����%�ܡ�?y򤪿��b~�iE�6���ړ'OV�
��e��br0��]�Vܻw���`��[�*�L8������U	��^\��K��9�)r��޽���c�&��r���%�2�� t�pV���_��l)�6oЉkq�s�[�PY>%�[m䛕��j��dl�'I��q�7o�>�\��6mJ��X#�� ���ӊ�J[T%��,0�Rr���4?���ϭ�7�	��ғ�l�,�����d�XWqՍBP�XR�cŉo�n�|�5����1X{\��-��QXs\�RW)v�e�q��m^Z_ $Vm`�p�%����k�/�Fћ �k�q�`u�F�u���r@e��ǔ��]�v��
T�"���Jl�r�����b��TM��+7d,w_�8�Ǽ����7��,�S�N�Z�T,�3��������51��ɳ�jŪ幐P���L��x�bZd |�f��p�LUS1�ē��O���e,11k	�KAfe�	b���L~�A �&6����V�G)��U��V�۠ĸ
�֋J��%��Ӓb�o	'$n���f�F��A� 6�#�C��ݽ7���gr�b����^�Bw̑|��-��&K���"��t�1o{�Tl�[n0
x}�1�R����c��h�"d��W,*�$���v�ڕ61и�� τ�F�"��)V�>�m�s�����M�k��8�n���kUW܀2��R�Y9JVq_�D1xՁnԵCX�,���ښ�u&`I�VAK�0��cV}���~i������Q��Q �h�)�U"Q�9�����&0�&1�*Z��L�߼D�O��L�P������=���`�"ra?X޷mۖ�̱" ,6Y��Ɏ;R�-�B{�; E,���(��B��#�&&�+���4�؝���]���2�������͸ۨ|)ic`��2��^���~W�?{nS;�ʭ�BH��TYPZ��K�*�W�1���"Zs��cv��l�D��( � 5���}�v�`0�[�%V �;�yMs�r;r�H�� .�ug�5k�$#��Sbe�_������q���*˪6/}�̐�� ��r�}�~k    IEND�B`�PK   �rZ�1.:�  )  /   images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.png�yeO�-�Bq����.Z(�����-,V(��Rdqw�Xq�w�E�J��H����yor��͝��I�L2�|��d��5U�	100��0%����?t���	��h�#7��'S��s�A_�?��K��K���������ח��孧���-���}�4��-p%}��c�4s�����ݹ��'N�"Ł�`my�׊��Da_����sY��]��`�~!�6F��	q�8�1"&��^��.=U��>������6�^�>1Z���� �Uw���I��1�vd�6ǐm�O�w�#T�7�<Bħ�O�Y�5��/l�8��)��*�ǥ����K���f�G�Dn,*��:��֘�ݜ���oN�`���쪰� �<)UjJ+��-ݞ=�T嬞o����B����0��p�W�	RC��r��",�¦��e��7���P�A�H�1��y�P,�F(�1}O���6ez�>�uby~���I��ڷ3��j��$<�洀H��%��;ϖ�o�V���$�=�+6��� �0����@s�	h'/?4�M�ίC݌ҕSp�u�~���-���x��귾3kF�&�>9�ڭa#|gTLw�ܟl�5�aI_z�߆f�~[%tQ5 ��:5���FjH��������fQU���Sז���_�8�w�:+ ��/ʦ+n�q��n��<�"��Ԑ~|���:�4�1=�ݡ�/'��^�E��8�t�f�x;;|*��ǌL����������4��?Ż)*�9�/��W���/.}�i�d͜���Ss72�6`I��3�������h������پ��I0�R��)#dg2�w �BP�p�N��	�
2�6�R�h���[��[�@�X��(��
O� ��A�޸�������A�m�	�Pn�*E�'��CC*c۱~1Қ"Y���k
�臨�RyL"W�x�E^��x\o�<>�|�z3 Is��$�[�I����*e�m�ȓX �рH)4oD��d
�X��/"d����h��q��}_W. �4H�$�H��E��k!+�k��~��x*{���Ģ��-���( ��h��(�|��7X]D��L��oۜ"I;ZCo
w���;��-kv�5���ID�Z�'䃨#z��[_IY .����S<_����cO[��u��^D����T�yc'�n��N��Y�C�h�ؓ��T��Ҳ���6-~�|j�������\����4�L��%-Q��ٔ�VZz�6��U�N��%Ď"j��\��!����u��I�l_�Q���w|{V��Ⱥ>��Š�����n3|x|��w��r2,p����m�W��s�I)�C��;���T���p��P�g8=�G�렶d��(��|�T����-��iķ�\�d�/w?Q����6��#O�?���ˈZ����c�\֍P�}0��G��۶Yhol���TC��F�%r'��l֮��o�x_���_����GP{0/�Z��Ӭ|F�L@a�.��s���|�3;�٦9���u�%z2=�9���wD�Z~"u�Nk��1y���5wϠE K�<�zzzB*������+��SR~����	G� �yw<QiG莆�������ʭ4�K�{��u���j��Ѩ�ft����q��42>V��CVo�!n�B�����=��!���_ʕ�c��'6��~��f%�k���&@��R��a�5�e��XDo�{n�̀}�wǐ0d����̓ �P�:������jӊͮ�!�Uu�7�Ќ�^o�S����܀��eI�s��|7%r�TK�������K�du1\a;ֳO!�Fz`E�����ބ-�����Uv�����TƳ.��]ܮؖ��.v�bA��.jM�Ǯ���������.��<���2��{r��""��Y���&1Z����׍���u#��G������o��UE�;�~ʰT^���]2*-�J������h8~�����s��:��~�l�h7�Wg�%�`�	_��U��:A��!3:iZ�^T�)��ʴ8Kw4\-�/��~;��e+��1Z�9\�ap�pb��leaE�]7�@s}t����X���� �Cf献/�[��u��kF��[���i�e�`��aS	mH���F�;ўH,�Q}C>�{��gذ|,��Ŗ�`
9�Ӫ
:P6���%� �84�H4G�b�},V���h�Bg�\[��"���0� �o�פ;*��Qv������p��3w�����J�#�G'Xq�i����"����Y��7]���T��'+8�9�$_V�TN��&�|�g���5�a$3����ܷx�fo`��܉?O�j���n����S��+�^rA�n1�b^��U�"(X�$���5��q1SH�J���Ʉ��$K�Qq/���NG�O0�h:�}y�[�.&j� �+�ma��yr���5��З�(����WF�&x&�4��[@9�ɪ�tmF�	����9�E��~�L��$*���\d�o����齬��߶��9�V��@�V�����'yG'X�R��M;�ˆ���%>/�$�� cv���T>��~�I_��~Z�Pv�޳_g�d�
U�/e�p͇����3�s�c�*Mi�!R�ث�8Y�	�N��YSud���d��y[�l����/XJ�v�)��������ٔϾ�fs��a��$�g��5R�����?V��-p�b����3��z'*�~wWe��F���9����W�B�_ZL A�,R�B��,zֲ]y��^ԺR���Y�z���D�J0I�"CA�����0u�]lC��j�� �Kr^!�������Tڸ�8���ϰ $,S����W�k�ì$*�3��,�0檋�K������j��/��s{�É� �	*̓�[|����nM;����3�+��V��G����<�0��4Z0�:G��Ps�Na�:�`U�z��������,đr@(6cV����N�ئP��l��;SE�6}��F���}[UC���v��Y�?6�j��\8�jabU�3�AD�?/��s#���7N���B�Cr�C)=^� 3.�_����1�c�1�t�I�9�t.�`4��
���M&q5�ޞ^J�Z+��1t��8ii(os#�6�(�g�=ϲ^:��Zc�����O��q
S�����!C�*�]]&mQ���%?"_* C�E��#�
��J!�F�]#�L�-s� A��c�t1s�[vn��qۢ6�.�cڶ���7��~jJ��:z�6�A�?B)�լ��c���n�U��ceII-�t���Y#*������Kuv�:�x�<�S�h/\�C@�Ο��˝��9Z_ز"�o�� �Z��].�9�ɵ�/�W����"jQ-�0�+UOQw��8%�ERV�.EbM�J���b��[�AA�&�Xw���5�C����B{�"����R7���$c�R�13���?.�T hS��e٬H�e���̱�*��Ҥ0�D7��(TC_�K��&b�	����zX����>}C��}$c-Ag�H=gwٰz����4V��MRp��ޞ��B�������lyyb6d�`��I��E�d�K�q]p�d��$��U�H�L���D��� �MY���Z�����*��CN���J�[��5KK&�����Q.4���������Kk��U�t,m^}hg�p���^ϻ���Y�6-�ݓ2:N�i��{QK1�@C=�0z�Az�=�PL!´��G.~�:	@��*�{��r�d��%^)�����������/���Ո|�b�_�n�d�'%�%�|��_m��zKW�#�Cͨ��9����I8d�봍��rS9�ʚ<gX��a��z��+�Q��|�l�,+�����U���ƉP�B�Ix����uX��с桨�y�q)>M6[�d� _q02}����IV1��Z�YzVw�|*������\E9L�%|��&���OI^/���P��'�q�M)y���(o�F�����A�3�^(~n��3��¢�Mbt�Q�0��[{�	��@�8���Յ�^�e��5�>j���^�@iI����w�w͜jG�RB���,���qK�qK��_q3�c�	!=uoGi�,���EA4�kk��=ҢB�}R�e�\�ቀ�]��[b�������)�j���#�&�4.�uu-�!�-�T�2��i&ig��p����������	ҙ?VA�Y��^NcU(x��J��ѱ͏p��ص�sf:��3^~#�=2ܲI?���嬸d��xN,��ΤL@���rl��z� *�Pmq#����__7 ��H�B<j'r���I��m�H�3��\�hxi�[�q�ӗ@[,������%����b]�pvR��Q{��̜�޵뤗_2�)y��ѝ,km�R;D����2]�L��R������n�h�9|X�q��a|i�
�W"|6^p�[�Wȳ�븅�`<kN�Ә���?G5�^l��2O�V��]7	��0��m�:���PY���&�%	'j"��,3cj_Ns���+`qA0


M�z�ax�(�)Ƀ<g�5$�0,�t�<�1ֽ���lj(�`/#�g��}���	,�}���8F�&�b
UQ��!;�b�#b'���dV����@f�(���\���S����#h��O�:ݼ��a�XVR}i�һ\`��\`��D�m�K=���}�ITw5!��	���
~�n`()xz=s�3�.B�f�X�i�k�%P=�Ԋ)�jcɶ@��q>t�M}�K�/xW��Iuk�[90��o�A��dy0*�I
0�Ά���}3�?�O�V�m����|4(�e�OӖ.��-Ɨ�����<��ϱ�#E��x���i`C+�D��+൐��T�������1r �^NI�i&c�u	_����xi~��j�o�t�>�d�S��,%��Xd�z�7i���C�_�{���⢫tA@z�.�S�}4%Ь*,�{�4����Dȩ��L�I���%K��g�%q���w�y�_�c�{qʺ�L0n"/�����zt�/0nGt��d��G�=�x�%;9����=�б����&�}�+�m��s_�l�bV��S��;�r�9�.W�i�����F-;6uoN��I�l��i��~C�"�p8�C�� ��؎�הݮ���%���l���ܕ��1k�:�g����=���{������G͈ne���$�(���^�������q���[�N
���D�h*��(�#Oht�aq�|*�t4E9��mK��(T���]a����8���f'��)��z��������\�t)���'�����`05�t>���Mt�=8mx�U��&��@F�<�)�^|�8� ��w5�j'�=�M�w[�� ���&�⸥��n��Ǧn�!��~a����y�
/����'��ڑ�9dW�����2¾5��.�#�쪩͋�@Um���ZlK`v,�]�#�>�7�1�a�d'�#��F\1�c󱢙�5��i]) ^�8PHN�=�"�D1��ǥ����аf��_3I
�G�$"8�0%����������������[�!���8r�kB/��S5c@B�ND��|�X�2��v,����\�)a�]���d:0N�s����o��\��ʈ��Ҥ�!Iu؆Vs��*X�tq�֗}Ȩ\��a��n�ћ>�Vt�ye����w4�F�)����n��oW��y���V��D�e�(/N�#]`z'�`P��ec�����H�Ħt�����O�]��B:�S����I�a@)5�J�z�@�%��9���Y���\�+���)��M���
J
G��y\�Z1'�Xߌ;���T����yS8����:j�!0-a�H<8���f�$��i+ç�t���!>�A-��\���ϵ�� ;��3��4o�u�Iw9f���f�4"�h�m�$H!{�O�g�c��C�C�)��ঢ�S��"5<���3�o�9���fK�!.�������f�^M�Y���T&۴Js����n�"��B�|�o�[�9l`���2ˏ��WC5���-�Z�C���c�zo���=^t$�[&ˑ䨤}�JzgM집D珦=o�M�[N��p��2�u�kx���ڌ�Ȱ��y�+��.�T2-�SJt�-�k��]��.��0zX�h
��ڒs�%�E��>�e��;��ã�/fMۅ�]j$8� LA����F�TM	��{|��EWՅӀ��"�õ���y$6 N��jC�^�&^k�DL�Л鴯SD�i�yr�,?PC�b�^����N�y�P�tm���� w�~�/q㵏���&����Uq�б%@������� �U;��?oT�-�S��4�j����JX�/���yH��v��Iĥڰd}f�kه[�[eo~i6�y+[�2�Pw�2Md��7"a	L�I!$����GNqZ�m�8qI{���;Y��l]�u���������Yʖ+��_��y
�.�h��f7z�\U���}�S"�y,�fP�Q9���5XeYL��?�.�������]���+�Z��9�j���,�S��~���:�=��������t��P����E����@tuX{V8z?Ѕr���k����7����+9�����뢓oC��f,�QM����E�-��M}��r��$����:�v˝�G�4�]Bp)���q��-�o>�����*֏���ץ�R��-�rc\'���F<�"������\t �$m��@p$���]-8�	Ǜ�&����u56CӐ�Q�� o��j�}||}Lk�ů�H˓��W緽 �.z���l�p��drB�1-E�� �G���v#q�߆�[��׿_A����h@f {,��ӤB�0�B�+9@���ȉ����2%]<�Ǜ�9����ɤ�޻��
"+�s5��I���N�t�{+HI�~���Vr��� �D��v<;�n��S<�x�4�at(�B!�n�#��J;�������>�Z˔z���L���:s�	����8���8<4 /���q���>�5���^�P�1�C0˓��2o�y�����o�Q�,VfϞ�իwCR�{�ϐʃo��*�� N�Z�+'M.��mݏr�)����(u`�{�e�M��9|����/GD=/���BJ9��.���{�f���������(��5a�vx�&�V��<䒛4���I��6�K��e�/j�k�Z�s�2+u^�����Xf˻��{k���s��ZY|u�F z}R#��O�:�S_�E�����ho�lW�;�T:��z�K��і.� ����mjr�b��lT:�˒�:T����Q?�y_��_C���]�3�^�I��.�$t��@��K|>��+�%�;&`�1�έ��9�s�@�TN�_&C~ͪp�Z����
HwTS��L�Pq�0;m�i�4�w{,X��+�� ��$�uԡ��ۧ�~{�Y>	#E;�D�YUq�.%�[��E��S�V���R��n
��O��:t�m�D�6TѪh���lF�J�ُڇ��Ev󧟿�
���/�������\N��#�_ J�Za���/�J�κ��Ȕ��w�QI��dˢ������j�%a�dP&���GW��W5v����n$h'Z�r��Q����R�.W?�MW� �Y󜖱���A��S�_��%=x *;��f�eA��y��#&�}�>`�k<+�z&�x���AC2٩���}ŽQ}ָ`��{�T���+�:�Q���}+e��T?P���L�"t��	����-T���hf�[KzGd��Rʦ��7�Ü?��	dX`M�-V]z�#��k�����5�>C-C�PK   �rZ?S��� 2� /   images/99226213-8268-43da-ade8-d9d07cfcec9f.png�gP�Y�6�3�3
(���J�80�d$g��AR��!I�,y�$9i����LJ݄&������y���s��rW98���k�u�k]k�C���.�\B d2O�VA H���$��̓�_~u��Q#�7��+��w|��@�� ���f��
|󆋔�������DrX��8�<w4�pp�Hŉ� �2��架������ge8p����9~�����9~�����9~�����9����D�a �6a����s�?���s�?���s�?���s��W��
?���|���t�+�p�����q��ds���,�r3�A���7��vaj�(��%'�	�ψk���XRKj�^ی�����~��Gz�޼nq�"�s�lz�c��*'��B���G��*����'�t�����Ð����9~�����9~���Fy\G!�~���AN{�8�֤�M�,�-�U���0/��w�Dd�-�h/j�`��z���L��qe%eP�Td6�`�$!{+m��+�H�0/0�EV\&.1����2wV�6Rer��t��=	���n8X|��^�V����ϕ���-¯%> 6#�
{q�$-��6ﺴGDW`�3�O�5wr�~�;�VNYv���.�7N''kg���}��:�w4&vy
|�4;�k��:�[�$���L�Su��u�w�4���Yz�+�,$d1<�nە��f�=*�����o-;+�s߾k9�����#����0I3��\�#n�-�1�i2E�=�]KeS�g�~Q���z?K\���N}��N.'�M��x)~M�銶w�����2�-#�z!C�܁�����k�U�<K���5,Oz-�e"l�k�xͦ�ٻ��Ǐ�U2�+u�D��uLǭ?U����{3Go}�5$H��67�Ck�g0܆�����<�s���?H�&�����i��rJ=��k���p��ҁ�Ɇ߿Q!aYP+ڭ�ұc�����X�."ί�b��$��f�@�ى�a>�[O��w ��[� _7+�����~g�EG�+�}X��$�qf��q�VB�<��C�����B�o����Y�xj������g�bh����>�ޓ�̧NLPK���ߨq�nd�����B�[F,���O����o��)<�j3����J�-�}^3�S����q�o�'<}'�0M�F��`7�bqmwi���~3��քQ���dFK[XQ�����5����b&��-wd����^H8c�V�g=m$�,�l~��"\D������ӕ-��/Cny6�*�)�O�|�����8�??~ZK��ɳ����[rm�2�#i_j>���1wY��l�[8W.5���P��D#熆�L<������"����Q]��]s��蕄\�y"���;�˰��G�v$��T��Zۭ*H_ݥ��<�>�e�g���P~8FoY"4���i�ɚ
�29�
��g�'٘,�����%|�}��ݙ�F�k&�{ټ
/���\�.���� B�v�ώwt�m.���v���2Ln�E;�3&�e��Y�zDU0�GѷX��R�޺f�&�]0x�;S��>	,	M;R�v�-�)�Z?3����Q��Hs��H����
�y�٩3摝je��4���%{c��E�[::4j���T�/��~)0���o lC�{�݌$O�4{!0uUe���1c6�s��a]�Z�~{0�X�����,��M�4-�F���z����;�N<"O�?�4�q��|�ɗ��Z�+у���[��*�������^�Q7�~����w�㔭�S'����:�X�,�����������K�b/~0
آ����nXn��z><Sj*<�Ij���}{��J��⃖��.���C�\�r�J�l��2�|�-5��u�I�>6k:��y`޸?-3��׺8;K�{�H��d���A���G˝�����ȩ>�ZhO4�h!5n]b�ݫ���R�4�W<+�Ej��7i��BS9n��;xZ%�	?�8 s�<n�%̝oz���(��-��J��/��jX7Z�����(i �_N��Z�û����y�soձ1w�7������2UOZH�N�-�Z�G�(6���oEuE'�pu0�*�S?�=_B����"�/FW=����ټ�*x'D}�}�6�
�����u�:�j��:�lГH7���3Hk��?V{�X�pEn9p�-g1���a �������5��!S'�[ԗ��<`uy��mZ����ݣ�<n�LKǳb��c��`Y�4=�t��?�����>n�~=�-?�1	�/s`|��R���x�g��i[k�����h����__�J�U:ڀ�z�L܃��._{�(�%'^�� �N�c�e�ڔ>���©��3p�B;�,����L�:6h�z���"�Qy�*��hu7r+�Z���y�6��s���Rv����Մ��eܹn���Y�ۏ&�>��[M�L�T	8��J��q>�x�%�ɦ�lx;��ƙY� �ZR�pf�u=wR>�:	��l\�����������(����`!�x����s�Z5� _*�ȩ��@�a�=v�0]��0�-�7�;��ձ�i�&�6_���<�Ik+����>fͨ��ѵ�N0CBK��R��J���j�u�X�N����{���R�6��t����`�g	nK�3rT]ݝ��B��6�|1��`Ba����9Ob9o4Bz�5b�V>3�s� �8	�c{7?�� ύ�b��.�l�*_����N�6�~?y���nTy�/~�8,'i<#��Q�n)��������h��ܖ���7��}��c�:z{��$6N�����:���g7ŎU4���4�}	M�M��f�5�����S��+��pz�e�� 9��BEؑ��#�*@hL�N��o���M'���E�e��h��$����0!���d����}) n�+�~�D�is�=`x�� ���q��$ bƱb��4���/9�0��������`6�������e-w��俀��� Ä1Koc�r�o�v�T"5>������?v� @(zP,{��9�/Yw9f�k�:ͭ�V��H�}��9�Y�o9Z�t��=� ��q ���[}�0
)���|���� X�E�������ѵ������M���Av, +J�X�<>��zFk`jF!(o�ӻ�U_;�����6}�`�p�=�5��e��������؊w���ǡ�����&����'W�Yɚ�HI�:r�������������Իk�oR�k�[	lJXN(a݃���-�������_<V��(��Ow�f�b��g~���ٗ�޷o�h��j�����铆�R�+k���)E��0�GwU׫��<�ݹ���Yh���.Gu>gx��l/���u��j�$y��h�����S�gE D������i@�V,�(��8,=be)���]i_Q�˸��|�FO�������1��U\�>ơ6t,��<;]�i���C�&?z~>%f����V�_���x�f+�,�`�����A`%���Iك~�llZ(/4��\g*�}�~�a]#�1�IK�
�o�z��bAz����P���}ε��1IŠEUUt��1:���0�{Ӿb�=�N��@��[������^4�7r�?H8qpߺ�yZ������s����~�y.�~�y�h� ���!~�2���0�����a&P�so�!l�;qp5	�RPW�hN�>���Bad4ڴ�h4�%ho��r�Ǔ~�}��ܼA������~NGǉi�_x��	C�����  �n"���P��;�Y�th�ԉ����M�!s��y[�y� ��2ǬK���CKF�4�f���ɾ
/��Ryp�`���t���!3��z�{F�Q\�[o�h�(�A��&@�h�*��E����U\��Hvѫ��Qx��0W���z��7!��$t��2���,�mO�����xj�ǋ���p��q=��_��7j�
���S� b��o����@�[�_j��(o8Z�W1 ?"�4#��ɉ	�)�Y��E��<��f>͝�M(-���}����E]u����&�j>��b�}�h�`�r��*� ���~�
dG[���s����'{k�����hvPO��L��_����/z��O�	��wK�D0�P\R����=S*���Mx�vh1C�cܑ��U������z �
 ���Wx����ܽ��aGn�s
��P� �����@���Z1��{x���+.~0>�[ ���큖Ԝ�jWGwynˏYC���ì+��֎������<����jEmX^�J�����d!�kEE-��������A~QD8F���İw�&~�p.��B�� jͬx��� q��E2�@S���Z� q�1sv�t���+,m�@���l~�5{�R|��� U@|��40?��m������F�O��f���:���pi��+0G����$`�ׂ��g���Ϋ���>R�Y�U_���om�MT�xy���]��;=;+�� %Y0fqiCܱ�>A����V�<��P��3�7�mf��w����pg��j�@�i���a��R|�R�0����hh�2�����_w��f����������Oq
A�j�a{l��������}PB�~`w�>��&��(��R}þ�E����o�9�X m%�s+�F�����ڽ���%q`�y���S����9�$����i/F0U��g{���O=�٣�;�^a��SBR�pt�cݛ �d���[����ef9�KA�v
��\��|�̜$�JN��N~u|�k���\�6�d�/�1fTpxog�2���?���'0]��z_[hId�߯:K!\����%8����}|/��FV ��((�~��rV�ӓʏ�x1�A�ܪq�ַ��Ԕy����� J��R�eT��m�~�ǡl����D8��\ЃY���}����;9��}�rR�ܷRR	3ƒmͧ{��8� �(��*��XD��b��2K��z�
���ݵuK˃�)�Qî~ȩ�PNh���M�,)e4��+����gp�X.xtd"��U�gS�xmخ���%Ey����ۇ����ع�����)c@��r�?{�TlH���Fn�U8CFf���������!w��|#���(p�7�x�b��6�ii��}6����b��?tG��g�K�R3+�or� ?d�G^��2�e'}5��Yb���s��+�_������5��ܤDV9�P�ׯ����^�

��3��ׄ!Tφ@A{5�E]S_EP��GH�l��%��a�y� ��#���L��RT�-�X2$ز�L�ҧg��Z9m���D�\�J�+�rO�ijJ����I>-��y֕R��1�#��s��j�"�饻�FoP��9�*e�F��{}O&vd�ؖ���] ���<a�%'���FFJ|#(��\���-���XcU
�{m�.|�Fn��@���:`;��߂!�:�$��I��-����{�	�+BQ*%O{��N��d}��K	�����(��r�������}��`���6B'��rV�FYv�w-u��adх����ވ}F:&9"R?��@];�X���rb�SW��>��'h���Us��M6��i!Q��oS{9ʖ������?,rUPȴ_YK��Q�QZ�����ҽ��d�cc	2��]�ZZ*		�q��^�k#>�xlE'�
��TyN�����_�?[U�ЄL|�ܷ�����Рd��1C�^�J ��8�(#77��W��1�G�`"H�^os�>������_M}WW!�ӗ�֫���Q��1�Y�gUl9�_=$Z�,�XJ���Bh�>P7hM�$)~JF&=��(���`=���ֈN2��8:8`���_�v�xˁ���]RD�;;;�����bL8ʇ���^�N��[X�����d\�DaC#�:Ϝ����Z_��{t�w���I`u.@f�9J���Q�jk�?G[�܃�»�49]�����­��Nc��FCO�]��I A0�N;i<����KV6k�$��%�.�<���:��==������*��pGx\-�w��G��v�fE�#%2TTb�����7������A1M������ڊ�ܗPE���͈]?�'��B��hg_{ܓ67��V6��/߃\^��� >��zm�D9�̮]Y�3K������?f�f��9Ɠ��-��M~g���_5�l-#� 4���lA��ʸհdc�m2��h��"��ۛ�)�j������z)<�>'��)��K�anD	U�_A�g5�!8W �F	g���'MZM�vy��@���5"���9I�/0�;ux۬�.����A�N�*Ha��46�M��<90�QZ���_��k����y��mv
MoO��t��ׯ�+�˼?R���w7&&���\��}W��2�
�E
�I�Y���zC�Vq8�VO��z:III�+/��v���|y�}�.�2(u�٭[�~:L<�R��%��5����$�&�f d�@}����A�q���~��a"��b߬f�+K�U��S��t"��LU���Ch����2Y����:xP7�op��ܑ����?��k���$~6RH|(v3��7�~��s����0u��8D�T�M�Q=��7����}����ct��is����F�\��h�_xG�u�<07W&+�H 6�ZI9T�V[-��8��kO���"@��(�LN=���C3zCqPgHb�+)1�\�輏����}�>��v��0~ܚK
rzg��%%>�f7*2==�i�N�8\��5���?;M0���Wa�B�_u_M�/Xgm{�^]���<�<���ֻy��綩.�g-��R����oH����? � 4����j�I�l�����8���1����m�\T�q>�gk�01-1[����������z��%(����s^�d}�<=�����8`��XPK)��O�GEP�,�A���/��mis��;���k#=��E/�]lJMO�̮�0��m(�uA��:%���;��I��o=��0Fo����7��������� @�t��Vx�,��g&����<��.d���yVOSRn�Jk))�'�cHS�{�r����u��&[�{=���3WI��.�`D񵋬 p��'']��WM���kyz!n-|��E���^�sJ�X��.%���NP6�h-c�(���$mm�qY���ujj�е�������1f.i �[ix������N���1	�����v�w�c\GO���0̟w�)rߙ���W8�M�������:)�q��- �s ÈL��V�?J[��Ɛ-��蘘��'u�ZxV�1���c�Ų��t���3�e9�J��� ���*k�,���pt���:�
h#,|�v�r�[[3$qq�]��}��\�n����oԋ�pT�A�対��]�f�5A,&"�a`>S�!������x�!��w�uX�&�@vq��5sߠ=v|��� "l��q|_�[�?^�Tt�1fخ��K���Jyh�@$����<
��,|ji}�������F�`�^⯰��w������H�A1tt�+}c?V��Q?��'px7X�5ޕ�h�o��DN2~�8��2%%4��������f�A����i�!(��
u $��SR��tt|�����C�!�Z@/�o+�{�i���hbR&'�(
�e��қ�1�̋\S��$9#J���*�:��P�J�P��\�h��\�2�u�Jaa^lT�.�p�a�� )���f4����W��ǝ�� L���ό�z� ˤM`rI�?o�XWg��}����Ȕ���"��'�3��VT�kZzh�Ǟ�.ZP,�_��U�ЧOd2Y_�C���jh�f���z��!䏆�}�nI������P�#Z{(c���������b0�@�bv{go�8?��~DD�ݾ�Bx�,ϴS]\�_�M7�w)Bk�MV������=>	�����ק���6)�q����o�����v{�Lg'����Xk�
�����?�ne8��M�K�n��Dw&9"�LBK�2Bc1;�ާ���ʐ��3t0ם�B��n@e�**`�RS<�A<o��$�����1����W�I;��V�_�pp�((�ο{�A�w�6B&���ق���V�����*�Бf�]w���♹�0���V��f��jN��:�z��Ʉ�Z��m��l<���_���X�^���ʰ�o�Txl�Vj�-`���xg��ηe��8�����m]�@���6�_����Ԕ>lb���mH�hV[�44���Ԅ�)R�y���L7�܂��(�w�A��bP�T��b[*^dL��+烲��ꊠ���̟\���C�&&W��RdL��Í��0�F��uV]{9 �^V�~~-��E:�
Sz\]N�G3D}�,�jkڬ���Z�?qssu����0{j�(e.N�����a�`�+?���:�R��cN�����g���,~���FQ8�io%G����u9��F8�h9����е��Y�t��qպ
5��c5���S��oߐ�a��J'>�i��Q��jZ{�"&�j,����|�������@g�����K��%����$PZ��lE��Q��O��M�`�(�����11���}��4�V��0�x �s?jC~�E���*�@tԙާJX� Xu�:��=�:���΍��X&���s_nnL�R>�XB�,~�r��Iw-�����O$�6�h�ր��Q��F�皺�)�}�ߟ���������-Q?yr�P���X���51��Мm�u��#ynh�V�Ųk���c͆៌���4���x&��Dz0�G⳰��q��I]]�T��F%� (��N׷Dh�hB��<����h����\

�)OQ�s��������LK�ӣ��p/pL�&�U��V]�m�� ��a�� �S4M�[˓��4��8KT*�4g�U�=��s+&*�Ã-6Z����6mw��(����Oc��n��89y��'$AN��������7q���;��T� #��c����V�/ϟ3�3>h���Ş���#7�{+���_��� ,rjKv�wP8�_jjR��kI���K C���I��z��Z(��wuq�gap��G$-A�I��c���śx���@��׵u��Ζ�^%8)o�K�L��`�z"#O}��Go��)\�li�[�����Y
��Xik��JFn��--7�5����E��pt��]_w�Q�~NT�^)�w�'��؄K�� b��h��j]���͖0���=��Hv9���K6a��k�K����4�j��JKҪ,����eg����s�y�����Ѡ;�ɨ�'�z�i�x����0nϛ��b!�l���-m/�.���D��2CBs'X#�X��;���p�Ç����BIC�9kXY���˝z�M�JI�xQv��D����5�T�[IA�%:���B�l�A�F����A]!�zNR71���R�������z��*M�.O_��Ћ@��im5������h�jg�e
?6f�5�Ɓ�m��������}�$��#�r�Jˎk�]_~����WRD��g{��wvFs���㷁 �|��!mk��/���0Җ��q"��E��G�3�Jx8n�+��_�N�uaH�4��ڕi/�[0�T��&A�S� �0�GR2S�܂bKE�6�t�~=j�%P�90+Kek��tHH��"qyy�.n�K'��YpG�F�b"@ߊ߸y�#��{=�k,�']E�ȴPe���"�������h+�.���"q8�-�7n�fXXZ_��y"mHZ+�����L��vF�5g{�Q)�ʤK67?�%���%(9�i��?/�B������3���А
R��S��)#�����m�^\҅|9�X�{_�P[�ۉӒ��Z|�U5w=�1l|0;����/W�c>؞�-M����7*"n�M��h�T�1�,.r2r��/�X�Ud?*)��P��S��'  ����~��e4ZI�e�������h����sIL�5@1�y�p��6��l�;�K��ixu7���߉t�*,tbz,�D�d/]A�n��&Y��\��\��)G�e��Eʏ�2V��c[�U]�����ڭG-�,(ߺ�D}��,�"�2+�����BMM�x۱͗@oM�		�ٯ`�����-�IK;i25�_����;�(_��u�f�dѵB81u;������p�CY��9jN­wH��1 Z���|Z�O��@�L
��q��x(4����h�p���,"qgU���u ��9��h��~`g?�T[ۜ5�P��< ���/���d�*�u˿C���?��gW����^��q/����\9��HJG�;��ejlx�		0DF2X\�p��Z4�e��
��Ϯ�L�_bT4� �h�$��l9�X�*�B��И�
*�Е�į�8�fnvvН�Cz�-=lI$���dm����{�e��M�
�M#f�k��X��p�z�x/�u.8g�
�����AIO!)��T�č�Zff��y'��܁D'�x⋲���iQZ^u����������sq�	�Ѕ�v|�wr���M0r;�(��}�����z�:K|Hp%k�[� �;q�|�1�>.]\�$4t|תʲַBSh�vXL���b��Ћ���\ˊJ<��
M�ſ-����>��3	ڞϩne&�������i>ܛ$>CfP��d�_��Q���Z@�s�?�����Dc*F�[k�.\�{hx7���u��:�l�+����i0�qK���(���v�3�4W���N�I
�M����]]�=�M��"�`ՙ���b<^�86F���j�*��r�N�Ec^;�����(���Տ]����<�#Ǒ��;���n�&2j��V�5gKc��Á�(̇�[t���T7���2F`.d�/���ė�O�a�	1j��>�L�}s6�mss��F|����i���Q��1r�( >����g��鍉/�'.�;T������2`ND��)�(�eF~(4T��L/?YHIq��p�6Y'W��$�{]���ϯ��`�#G�Ǎx���2�m��!��~�9�r��҆�թ�MFɬ/P�i�����bԨ Uj**�����_u}��ыJ����>F�4{�)9}��P����4����ќ:�����X#�]1�CR�wa�UW�-z;3����|"i@_��DI���Xr��B��U�B��.����;�z�;��A~�ݷK��%i�6���T8�����:X��x�=��4�i��Q?�Bݬ|�>�@��h���֭3ۆ�/�i�ߦ�_�>hR�H��'>�W��XK˛k�ܮ��ZZ����������X�5��2�k�vq�$b�e�"Ū��l��PUG{c��l�k�Cӊ {� ��n�4J(*L�vu;�^�G���Zd�" 8.9x��V���FD�C-���j�C�@&��l��J�M*+5��k�9�i�.�e<�!QQe��;C�h}ԉX^/�E��ep��E)��G~�j�n��j6�����O}̎��San�q����O�$�
(o6#.zz�����bNX��[���M�l�ll�@���s|i|ӑ
E<kKZS�M��ׄ��<36�[�O \�Lf�X�h����_C�_���X&��,��ǒ�.�FƛOa���a�{�OU1/���7�@{x�OSAM�Q��w`�����5�k�AA�J������>!�4�qF7��$� ���t
Ž����)�_�� �܃+k�q�='��R4�kr���	^m��[5�,
�|��3/��#�E��wI8表~��1���.�(�'67���
�}v+#�J��S��Ђ��0��z����T��g	�\��?���{��x;��V@g*��1���`�dC��k3�J���CG�$a�'�Z]�����Eig��P�>JRP~������.��QM���|��fa@��Ȼ>^Y�6����� a�&'�����[���p[��"�Q�7+{�ui�kC�|6袵��Lm1��P�⶗e섆׸Y%��* !_D0���/�oZZ� ��]N���Jq�e�Ǹ�k����Zi��b|���:;-/�O����������]�^����DA��?�V�����d~~q���¢�t;R�-�`��%y����QH���.�qʌ���6�鋵.3EG%^��c���$������O%$,^�1�!
�T"x/ܟ��ΞYT����; '��hJ���#%�8�]@�G�j0��82�+%2��U����h�˴�@>L�lĠ��m�0��T���B�}�6�ݕ��@����ԙ�k���m!r2$��������k��0:L�B�����A&`t��sV���l7 .�_��*��"I�+M���N����&j~��ϫ+CT	V�����F	BN	�@8��S0N��)���<�h?	`��[ b@x�>,����_=���	v�1x��e&���k�}�_Y^�b p�*�g}l����y������,@zl�9p���D�'&�$�&	;�gxه����:��NWAD^��!��wMG�Ga���̇�x2��K��X�f�� "ˣ ii��[�-O�M,pB�e��F+ˋ���Ê
�����P$5��N�v�U:U�['�}ț@��e�����+\Ζ��wL><j��A����tt�A �<��<��6��a#}�۬�3(�-+�ҷ������kkׄ��)�O�lA��NMk&�͓\���L%H��k���=9��u��O]YQH��ڠ��d=�%b�a��r8��(�N2<u�\n��J�{���� ���`W�Mn![:<��^�IlW��w`�'��ޏf�wu�^�g�0�w���(�3:���p�iy07�	��Z5CO+��^C��("�7������DS�:	�Q�Z=n���$l����E0�(lʰ�44����P���-k|�v/ņ��Z��)��Cl���f	�!:-ϒ�}ך�����m��M.�׀vJ���V� �g��������O��I�t��cq��\�fIHI�q�����-I�c�#��4�4v@�_�+*��A'z���fK<�k�a�{.)�N.�0S��1iP������@��<��Z��u"�pӧXX'Z�e���,$�]q�L�Rݥ�V�u��[7[`I�\i}��#��$FF2��\���K�`����N��xp*.*��w7����?}"]�0��X8�+�{�t�<{�,F�t`��l]Mʳ��?��Dm������M�<�
֮h�<��>���_R$G;}<�َ�ш~M'���}���}yAi�,׊FBw�I�̣��e��O
��VL�m��Q�����'-~dS�N��t��uOο
��j���r!�	���t'�7�}N]�GU�����o�7��mnZ�W�����2���3���%���ʭ[��s����L@�h�)��͌��[�>�O^�1�!��AI`�9!��d _�[��V�s��_'ײp`,gc�礯/,�kğ7d�=�%���OC�K�����蕾�$���w��sUnѰ�{�S�)ނ}�x����8j��|�;���a,)�m�m����I)�=1X��N��������%�=�5�<�B'�b𣞫 �*����H�
6l���G����#��8�Y�x��h���9MQ�Q �D'�Q�~R��?�ctW�b^v }	k�9����Çɾ���{J���A'�G������|J�y'w������W�_贮��(h����`g	)(��.���
ߏ�Y[.�v�����	��~4���$%K��ߡ���y�,
�k�/�ΩU��ԍ���-�MA��gB�U ��*���
�Z[�$����*z�	���g��������@d!�s:�9J�Xٛ�����R#�S"@S���E_�n��+��NH\Gt3���z��ʧL��r��q�Qt� zj�u�=�:�&�6|��f�J�֑��(��{��PuM�w�ѯ2�(��8s�W�py��	�$	�ߴ>��Z�b��Ǹ��*@z<*�����rr����x�^7t��<��Q�}�/��)��o����]�q[�7Wl�����Z/{
���F��{��[_J��>  �#�N�%$����C�#��*JI5�/�w�K³���;	��mp~��#H�If�꿠���P���|��4�TUf�'@�T�mI�3|���(��Gu�������4Y��7�����&0H'�n����H�]Mqz��,
���Q�IuQ��@,�C,V�e��W���JȾTT=�b��@� �FQ�};�����Zd������Kqv��-L��$}�w���2V��_���4/{�aRC��xYZ��X�%�q����J�ͳ�!1GM���K�*F��I��;Y���2�i)N"����둯9`�g�݃/-f{�T�}�����hj��U)Wע�JK�lN��ᗾ5m��A�)x+�#[ڏ�����#���5٠'�����_�9Վ3>x����O`()5X^��t�g~E=��s��l��p[�"y��Hk�4������B�]�0R�}$~|L��  ���~�~����4w�)�Xָ=�Va�!�^^��#���}дG`.ɔ0zlu���ǿ('�m���3m����D���f1�7?t�T� ��i/M Q�ꞝu-h� �Z���\�,��a��M����u�8��i�pt���Xt�ũ�J��5�nA~s�:+�_f��!���l��� �Y�I�\���.�,�z�ɪ�����o��d��;2´"�ߌ%P��{���IlR�!���<k:8���XE����4�~!]�g���5��yd�L%�����-��]��w�{��(g��_2�U�e���E����~t�קaa�}Z��/2����v�W�g�Pńw��x�{X��Tw�{�@�U3_%]���$�j���9���_a���\�UAM��ў�!h�O��1�"�C�g��|=�{/	s%O��/�U���������XŤ=�����.���4�4�VR-���h�%� ��+˜�&��;��^�Wx�L>�e��Q�5<vH�fB,] �����;t�a<���P�R�*��z���C�(^��89���8�(B[�	?�C�zY�o
��=/c�"t�?�t�+[����ɲ���>�2��|��I��r��;N��{(}���|м�0yeC����n�%h7�!�dkLn!�%N�Z�	aL��,���EB��Wmu'䒄�Sx��M]>��g�g�NN����� P��������ꊕ���ԏ��H-�����fろL��E�=΍���p'�i�H�VR�������T��'wsN��7���٧�DA��%�������@Cq"��İ�YQ���� �=ݙ�e[�Ԩ�7]ب(ttQ�nH��LJޟu���Xzf�~@0��.��I?Z�}��ӭ!��Β#B����޵�t	�j��Bt��>�W�����Ԓp6�x�8�Z3����7H�\��c.�&J����,�Qh겳׮�D,v���u�O�$�6�����$z����={v��*��א��	h��$�w�f �t��,��_����ٍp�ٟc�K��L��0vp��T�. N+���m�]�{� ���m�'���q�h^�.:��/F�k�!_9�)"�I���H�J��ϟ_2�:l����o� �/^��^i���;1�j�>�=��6�K�Dr�.$0>m���;�	,6��<2;??�Ț�!���׷�͸�o�����;l������x�����㳝#�\ۏ��S�����^��R��>�L�nj��#ܜ�:�?-h-���)a��v&\���K[ŞJ���O���xɀ%�Z��?���cw�X�|�4��O�4�vh:��EUS
�zϵ����
4�{�X����������� @�S�`�)Ǹh&�z�.�����O��Ӝ`�l�FL���i2�Ny���y��F�21��Z{׌��㨕�Ќ�i��˵�ҙ�".���e��E�(�]\��@��+ ��\�T�RxKk�+�#�dZ�+k�<}���p���%)t�)���P��g|��#���	���ieg���O�+�`&�[k�*)�Vgd�k���w��|~OD�w��5��n����5�OP6 N~#���K�(���3���/R���.k�juI"����8Y��.��C�ss�����ș��2�J��	.�a|��;#B��m����B���dL��u<6�wK�z�yHē�*�&��L�����~o=y͕ܸ������x��~�Z`�Pp�o%��V��%�~8�Нm�[4\h-��kp�*�9���ص60�����闱��G8�aDD %�[���Z���(Ι���s>��y��+�.�����(q˯��oEv��d�]��(w/���{��{>��9�+@��tgK�9mX��ɞ�e��ޟ�/�{�O��|v��q��Y�9��nm�\~�{"���)"���|nO>?<��vz�����*�M�z��X�ޏs�݊�ޠ���@��gy��I8Ԥ�*_Z��Nl��y𜻢��g��Hj�(7C��x���&p�b�M�no�i&�Qi[�g@�/��0+8�qh��dٚ70�~~���p��+]����]�>�,	�\++�Rj���Yߞ�c�4���n�����f�8׶H��������Kw�.gYVWq��<2p��3��^v��K<�����|���C0�{$NZ_���$Tq���{I�@����ڬ���%/��@k��&j0�ss����5h5�ݴ��Ao�͹�ϙbQ�Jt��wF\�b��7��DӅ�!��`�R�fg�m���>��+����a፝��̸d����;�a��K>̅V�����ӣ2MT*�{	Y�����Y	��W���@<�cC���[ݎ��V��w�;���9b��
�E�%i��/��s��i�~oRW3�+�[�ML2�w���{���#̖��д���д=ר� �E��NDu�sV���ϪF�)~�_w��>����nH��>:&I@�$FG�UuC|��!J0���@����GS�o.\�鿨�h�Tij��{��F_���+BA���2��}!��U3��2}���_&�^�.:R��;9���i��L ��=;%e}�n�K*�{�ueŝ��΃e�:�ϕ��ؔi���d{{{U�77��@�'��{�B��ZU��Z��T�*iE����B���{Qt�l�]-L\�R?�a��<?�ɾ�b��s>����~`n�2_���-����y�(ߔ���6I�Ͷ"�i�+.qpH���A�!d�U� 1q�ư����qO`ڛ���B�9�z������N���[���/7�+���иDv�!e� �|�x���+�j��_g�̸z�;���xn6�@W��^�@�Add�a�u�"���2⿸n��!�%�c�0����,�]���^�T�I�T�`֏���)�\��@z싈L��6=�-��H�<wmm]�-�����O���x��֖薨��'XAԻ����-��'�s/��<�dC裹g�g�v��'�
Y22/�ڻ�<=�
��J?7�����w~k%O��77�Y��y�S��ŵ|�{��g��9�WQ1@!���}����"7\\�������CsN�CsJ�w�H�&;@v��J��x �1%dc[l�2��g�Nb�&�!��2�#&t���R���V�'�ÎC��v��� �U��Q�Q�뇱�����}N8�����¨(��?�L��J{��dS����F�^�+XbH5S��R��V�H^bJ�Y��/�a\ŧ�l�A�\�w�	�P��z�O�A,�K1����2���F"H4��.�D!�5r��,'�}X~W�ʜ7�r����ωJv�Ƣã��y&�Q��g���ggA��
 ����I6%v=Bpm$h(�~F��"pc��ɧ����VB�=���y�4R�d&#~�"UX�8�ʃ8a�&�T�ʺ}�</x!ax�,��-���@�YTb9�t���U ���;�����r	�^DIADE:E�KP��[)��V��ne�ai�.�����g����8<��33�}�=��y�O�|��,�k'	���P�T���{f���ec�{�ʏHD��*�/��X\��uH�%���ү^���Yȕ;��G�3��R���j�=sPr�B�]�{泛S����
��<+�$�����^���F���O��4�Ź�&C�\1���с����Ξ�O��m+Xl�����(�:��ڝ�GW���.Pvo��yR��p5'��:b�_Y�@O*p��Du��Nt1��"ՙXP���f�'��p�bvy��EF�D�*����w�?����!Z����!�̽�e5�h�z���&T�]���R��ThLR�9�X 7�����l�����NC/nq�i!�u�O,K�K�+�urf��vk81�ʄO־���#�Q��ږ��9�u�0�X�s�]NW�y���U�p���rIx%�b�	�\�B`� �E��ilS���H��Lޤ]<����h)�kf��?���<�e:@��U�紜���u��:�����7ׇ����.	��?^�r������c�G�۳Y�[��Im	j�c�Mv_���k��iV�HP����v����_�:Z�';�����L��=�C�v,�D�`�����`.�PR�h)+IzY#��p���|ՙ/�1`�bl���՞��rX��<
�xJ���וH�r9�@
�9��Z��-�X��6���i��mP���Ik�D}�]�onu��AU�X���^��S`�{R�n��<�澁��R�7a}���~�+a��k��!�v��1*_�vKn�T��>d7���Tn�}sbA,�%yj��T�!�`sݖ.c��nL2t�w`ʢ/�F��#f8,A����n���=j��z(.��v���:�J�͆rqm�V�� R�;6���他�
��Գ�_�����v�N�\
���$�[��h��";���[V]>?�����1�J�N�?��/G�+��2��`��vw�+*":������w8�y2����zh]'�nWex�Ӂ�s�o��"�-A�%�jC���
]�x:D�2ER��^;�Y%������Y�8)w�ʷ w1=�W�������W7�b��`��Wx�b�vw��_����$�V�*�=H���>dp�3n^ǎ��������xNg֍]Ѩ6,��G=��XM�g�|�@R`�&�#�������*|i��%��P1��P:�0�̧�VC8d}_����%w/o.�}��6�\��"h:X=�_B�6�4#H�b��x֡�!��$�p=S�<�QC�А\��>翻 ��R^�sv�A��{��C����c����R;�����Nj�&̐wpwޙ+���o{�5��$�e��:��qK�9o�8�L�'_rC�|?teJ=1R}[�\�QE�f�7?�j9���V���AJ�ȝ�Ro�T`]��D[�uĖ��Ỹ�����(uv�7�'��-�w[Ìg�*��L��A~�L23#p�����ٛ�:�$!#�Q�t���f>�P�ce���:n�R��uH�Ҩi�M#-�)?�_a���3>��r�.����$�н���3�y��F��$p+]Q:E��	�_��6�^h2Y������B��
�f��S�O=��%�v��T�.�����l,�'������M0�͕n�^�&pX���[ ��
�eʿ�`%���ҥxJ3u�֏���+�R�I\�߆2�bѹqDn�܃G��~����S�p��#���jSH��>N .T��+������~��?�U���Zæ�X��HI"`-�?ɐ��XHov��i�"���AoT����UЩĬcUSw�+Y ��q���eN�� )E2R{���ϟ���gu�_��\h~�(��(n/<�:��Q}����� oԕ���^iW�_���)��S���=�>A SR��ʼO�r�0�?���+ʚ��ߺJ��n7�oq <+PU�P�,cN%b,�*��\�8��ܜ!_��l�µ������<��;�l�����c��_���V��y:�$�^�ٟ���`�(?�n����9>9��6����k@A�SjkJKk��\�MsYX&c �&�+�Rb3S����ŭ�}W@�g����R�#�����	4��87��W�8�i�"�.�ꁇ���V�����-U�>XP���/)9c��x���U�:��r/�>�}ZU�v����h�Z���a`��Z��Y卺���c�W����acK��Xp����6�Ԕ����n�H��U�',>��7�nni�i7s)�ھ=pK�Ǯ�x�wdm��~v�}j@y�����cƨ���NsC�껼�D0�sڕ�V���}��b�)�[�L�])�FH2�w����2MȪ��>|W�� h)�h�?ɬ�c�
K׿	S�G�bAA�4�@Vf��.s�^��w��C=O�<t.M����9�-��fG##E�����V��V��-zn5f����MZeE���d������X�]���l�H�+�$|q+�Y�!oS5�GE�yr��x����G�kD/����M��yv{j�uu}�;�&e}R㒦���lf��=\{�g;U2����M*�.ì-�_�%#����u/N���6ܘ��!�	`=��>���?�(rm�j=g� |o�
sq��\@ѨUځ�1|7�����O�]�bN�?�Z���,�T�$a+JQ��{D�Sw�b{Np�D[be������^<�ff�}^wE�_!2�$JKH>V.<���݁�'����� ���0WP<�xo��U�9V�l !��j�VE�����	�:�~JV���a���8s��_�|�tg~f�1%�.�θ\<f��r��B�#�_�`_���*��7F�#JJ"�"?IJ�&��zIAu�Vz`����yHXϔ[�A��ʕ�=���K���hA�"�2$����mO��]V��[�y,����~1Xvp��ZJO���P�I�j�?՛���~���qh0�]�vv�=7u���j��=�T��{:UfffeT}_]�:�HV����:�d��t�>���\A��I��	�xn�6��{��>I:Ï/��i��h��!�����6�#��w!_���8ި��,E��:��'n���
��k��-�3��9%�AJ^��,--��x9�i�1DcՐJ9Y�g�6���콳p����My"����p��v����ڵ�]�R'�E�s�у�3�jχd�/�ʒ	!�㉝jz5$İ��j��E}֟�󊮲3Q�k~�]6X��1�������lyg^hE`vN	�K,S(5�&Z`��p��k�����,Ht�颣��	�%�A�n�ey�\R�����s[��d�7M$/�9���qN��r�}������T�6������5��L��R����&`$�e��GP����И�:�kH�W�v���W���\�°�ܯ��q8-<e�_�"���ú�~_�������ڠ%����S���K������N�����n �������:_1��*�t�_�O��˟a�myn7�\|��@�$ �	
���4��9�Y�������acl�z闱��BC{�):z�_��Z\����șt���W��y�ya� t����#�|���R�4�]�҇^�O��g�ӽ^��`��"�AqK�U�T�຦��M�&��jF��c�}�6�g��u�~{C�'!!�b��?��� S\Hn ���K��]AFy�O{O��13��/x�~y�- d��+��<N�e�O2!Jܕ0�s��S����8�?���W�������~<��n����9c �4�J���q����p�)}���oyi�.�;b6p<���Og�9Z�O	B���>��֓3Ǳ	�
��|{�x�.���J�	��|�>=zqUf�Di��s������y������P�����Bd��nD([��x�)��γsx�R�*����BՍuT�\�^$�O}��"J�0 ��,x*Ͱ�������m������/�MG����cy�M[��J�Q.{+�-t��/ar�[����V+��"��L�e[2��h��
cVr���TY0�D=��Q�3ߚ����M��P�{�:l\ 7u$�V�����~70��Gs�W4o=qj���y����7����f�����1b��D���XTbd�T˩��Y0�[\��tB����C/�`��)�_�'0��d1%���I� �y�|��ı�EX�,�+��H�vu�=�7�rƑ�ii��y9Q5N�s���:�v�L�n ��7����4�f��(CƧ����v��i?�#�����Iۅ[(��9^[�_<� �{p��2�v�d�{��|�)�)����1��$Q�2rEV����@�C^G˷,\��]y(��m�����,�Wb�����w��ff^C�C�Fs�2d�F�
^$�\�++�Zδ<2@]����\2��0��¨+�Pj����F#4������*�ǃT���P1M5��>��eQwF#�]�P`��w0\�̬�&Es �O�������.��*j[p����������D�l�l5���R������4�D�ܲ�Ng�t`����/����<����ꥊ��;,D��������!J>�4����}�s�r�����l�;o2�MM�JA�ƉWe>O�H����-�1]���j�k�[3�ƽOGmq�#օ�2��+����ػ��СV�d"�������$O��@���V9�0 ;B�11	�f����ZWG��LE`a)��1�(}|܇����C��o�뫬���Q�p�/X� )��n�\�(Ri��:�=����f�~-�	�[j�Se�$��{WY�����ʻ�������z�v��`e���m7ƿڵ�.vx=�1L�r��@����vK�z$c!]*\�ݸ�j���щ."�ә�%�d�EQ�c���\n�W���j7$0�'$�~r�E�N**E����?aT?{�ۖ�,=ѝ+���ji���]?'������L���~��m�e0�����:�������� ͆����}'!]%:rM@�8j?R>����m$��~��4T�`�f����촄_�Y&�jj0�r�s��)UB�'5UKk>��iT/Z��>��1G�%Zq������!7~Y*dr�v<�%�	��O�wR�6�}��t,3��H��ٵ��УNH�zc�1��~�-30��[K����D�K�Y����c�)�Ƴ��iN�t\�&��B��K:(��������M�|,�_��3MDw?WK?�r>	�l�[�|h3mtL���v7�rѱ��0J�'7�hՌ���yd��2��[�}��*>���?Cg�Fg��{	
��Xo�#"��AR<�/7W*������j��� �3�)�~j�<X����)st��}��?O��N�Q{���`pi"����@M���/���آ��r+y�� �'n88��8������{tq�Q�L��`@�q��w>vf1wµSR������i�́��^����+1 !����U�k2J�V��� ����F�
�Ry�;Y�O11��v�_p%̿��*b\�;��A2KlSIme��6�������V�"�����+6��u�ȫ�Ulum0�'ǽ"��SS�~��)�r1�U�K~qd�˺���i��P=;Zp�x'&
~u�n���&|�
����QYw��7?�bLZ�[���Z��k�U���ANU���7?uV�t�?׾�؛�\U��£�Bub0}5������{Չ17W#�$��ibl�(���h7���1+�ۈ Z������c���?0�;!��6<�uu� ���Ɛ�GH����&��B�1ܟ�S���|�i˪v�x��6����	��dn軉sS��0�N�}�ÅI�,�,���b����i�!���� =�l�g
`�|ߋ���'���N+=ۋ�%�M�0(�M8m��4+�g�!%���N����i)7��Bk�h�W�n7�����jq�����+$�1��hL�����K}� �eU�!�Rp��6i(h����_��s��
t"2(J��������C�z��Ps�߰+}�wAJ'h16v<�n��Qا+�2�b��s����_���?sD�$dO���M�ڝ1����b�R�s�ׇ�%�.³Aj���W����X���V�7���#��]ó�h1팒s���x��W�\��8���pMM�ט�@ʄ���'��F��!��=X�@W#�\*�[z�iC��{��4�I���?b:�w�/n�!eE9��{����3����E�b�H��`-�+[^��Aly���չ�Fͱ�>�YJ-���(��F%��/:�dp��>�/ ��x+C�^i	���q]I"�9�B@?,�b�{����Xl���h���B���i�;b&����Y�J(+t�!����Q��J�Lzv%����Q��F ��]���$;(BO�Ř�q���yJ���FY~ ��T��s6�â��o�i7�f@~<[���c�>fwu�5��`�
��7�$���%;32*��DCuL^Du!Q�y�C*��W����P�E$����W[@�H�G(o��~����������	L���P0��b`��tH���]NG*ͨ)�^ڌ�����jH�A��z^�xu��&�aK������#�Q���Kx(�	k���x�u���T]'�v=��Z��=�DH2�����ю!��\6�}�Y��gDM��,�5^_w儾���d*�ۡ71��[���F�+��>��2��1z�V�.�'�t�2���,YԵ��BT�ʾ���f�?;Y]�^�-6]��p�'��Ƶ*8}T�����݄ZqSdi'N� Fql�i^��::Fʑ�}��t�{w����եW-�������nNz����G׀Y�,/+�n��e4�!?�eB]���Gi��4-��e�����3�~}�!��R����MM˂Yh�δOmIr�����-'1��
'��>��9�n��$nnjcMҿ�,�1:�
E�Ʀ�g���)r�\�����ec�j��n
((*�]���ϳ����G���9��,/�����j�t�j�rt������ͬ!�؊P��6�`G�gᣓ�P��Ĵ�y�'A��G(uqޖ���V��%9�2]�=��k��bu�5A�{H�]gwp������7�!#Tw�m;]<�� #D�Y�tB`J�6y�ܟx*.frd�Re���j֑޼6�]1}��3b��C��(/��ܼ�i���>їH�|$��yfq|�'��M�.��,�_fNM���?"$6R}
��9.��@\��=?����2�Fs;Pmj�023H�tv��`�}�������=���Ѽ�#�d��
2��ݾǏ�����?�M��s�!��bFjB�\��O�J�r�񣝣	�TDLfU	 R�r;I	]��t��F����_��n43#pp���<ݛ��BÅ���s�0	�\h�����~�L�LKН�^9y���'�gw���O�6� ��P�=��!Y���
t��9 #�}��s6G-�硰(&^ݫ|��{�sQ;�??�iv��귯��jT�{�����d�ٴ� 3������*�,������)C��kdEG��2$0:Y��\Kh}�a�3���5e�u<\�}�-�#%��)�1���M���Ѩ)ٛ%��"�Aj�~�0����۾�K�ٺ FH!}�`T�����T���L�9�G��|㪛��Bc��EF���|�I�\9����Go'O/;?u�7��>�#����� �D�������"G�B\X��:UK�����DU���_G�n5 �%��SqJ9�tb_ϙ?�����j���u�yX���gCE���M�:�;ɫK҆�ӹp�`��Ų�.��zL�? `�E��~�]���}�g��L7�i���JO'V�ȟ�-�L��h$rKCS��2kԡ�=d0���A����ht�J3j�~<��}�^Q��6�РP��yy����du:��BQ�">q�c%��Sn�t3�n
�@����Ё�z�T�""G
���dyu��I�:�Zna��c�a�b��I�2R�g�Ǩb��\\�ڳ���kS+�1٣���(��.�H����b�v����>u��ϝf���7Ǥ�p�<�BG!���M<�vO��NIɰ<mi��8����}�������W>�u��#3k!��3
�MZ�΀����8���<�a�Td��r 쭿uBr�!��奬�X�m����&�z�����&j�8����A����Ŗ���ezŬZ�}J�twG)����D���ҐŲ� �u+������̼������w%��| �b�	2<s:��D e���p
��5eܘ����!Jƕ�w���͗�>�U@��o��/4A�o2n�|y���P�6����0�z�����8�EeQx�P<1��~����[�g��b����a9�$j�n�ru-��=y��=��5Zu!�	7ξ�7�i��c���!DI�2�X�K�!�][s��w9ZT�(�ى�|�N#"/�2@�a�����P�Ú�Q+��it8Q��;R�#WN��Z�'�)� �	��B^M��O�vg�nIJ�h�Ҏ��#�	�7�]��?�q˚��q�5�!::��I��%srl}�����5h��0h���"���us@�*]"J�si�n��n�oM����u`
Sj'���f�~��h�q+��i�ٹ��l<�X,G�����u=��Jz��1���p��Rɏe#r�f��6��C���I�de=�v�2��U�E�������8�>�@0�-�b4Szo����Z���M0���_�Y4���ai47/M��T�cb���{o��#��D��guL�rۉ�YBDީ E�!P!'.�O�u�^�XLy*`x{R���?:��ۼ��7���1)RP��|(J_��Д[�kux�����tEEE���c@�<>�V2�+H��r����S�����ǒ�W�>�	_v3����+s�Ю�ANŝ眸a�)p*��H.v ���1�I���En�3�
�I������Oo�b�t�u<��\rW����0��V&����pd���[�ۨ��eSa��I��mU|�N7��!D��S��D�ff�,|]:P-� �ws�CR��lT���M��p���u���}��U��ڋ���3��D�������bP09M'Q�V�`�.~͆��'ׅ���B���^�U��(�8�}�3/�n�ʿ�!_Y��:����P�<��W�^��z����7�4���p�GU����	uvu�H=�H=��zbS���$ڶ�:7�é�Ԭ���آ�_�=���1n0ra��d4��z��F�"!.h�I�Χ������6�F݉�.vZ��<-B�{��'�Į���&;0��YoX��n��){��Jt���g�H;�W��@m�<m�R=8OS[�\Z�ȵ�,��j�g�c�O)�1ZS%7�+�>Q�˂p���ӳfoH����AA�xL�<,�m���.�B^�i��1ϒs��kOy�<�!._~8-����-gv���=u=L�~{i)�q)��F�����gVK��K~w�ܷӥ�-3������7�R���E~@~��g�y��N۾���B���<b6��,"�bk�'�C3�B�AY:>�#��w�Q�و�P�B�_4��qX?c7ư�)o��U|���|	��o���V�Z2�h<�?���U�D��o�va��?y�7P��_����W�x�^���q�װ� �:�֬��u��Nb&D��|�%�]�r�oENR9;��ȏ��߹�8�������1�,���	�{�oLy��|���Eb�Ϋn��%f'Sm�*O~_%���^DYu��Xy�)XHz���Aj~�(�h�q����~����0�v����2<xx|T���,!��)1�g�w\�L�G_G��`"`��[���*��h<"l�2j��pГ"=nNBt��>���SX>ɘQ.�U��HR������ގ�l���M��n����uԄ�b�� d�z��Sox�[~p=��*�0��z g��K�����/Ưr֐�_��a��_�)B	�-|�tq���i�����W��Xd[�Gw?���6*h�z��x4�(�݉g[���=duGr*U�?V�6>6�L�ݒ�����_ۣa���	X��n����V�̊R��l�5�+.c⿜6@�����ƙ��;��yC�^�-x��VC��WI�n˹��5%�\8E�V�?K=.��埏��>���$�� �ԛ������r�o�u[q5����O?���DM~�8�۴���=Q�,�u�$�{��H�i�:�9�����Tkn+�B�D:S��ϖ�ͺ�5
z>�W�E|���^�H�VK���1VFRϛQ]�*���-C�PX�^s�����B�t���iːV���;7^�6Dbt����/����#�Z*)b(�(�!H&nn.P��w�×�x����xSS�`�%�RS���I��P��оJ;���2��c�������E�+-���P֨��0�e�1�r��̮�^q��Œ{���_^���\;o�5����4�
rΈD�^<�j�V���[`�����җ鍍|u�t(�P���C�$g��q�k�qQ�)�`���G[��[��B�M^�Pp�DFy�{�����>�0�E������z�gޯL\���2�V˪���x���NK����S EQq����$�[<[X�m��tk�a6j,G�����S���b9Y\Ћ&�:��;kW�d5�;}��#%��,M��mr���11C����7[�/X/w���G���O��]�u�GX���W��:땓%��-��;9O�yAZ��#ڠ�@���8 ���q����Q�rλ�O8��Ū�v�+�2'�&u�pQ?�2]G�4%�*���>u_h�a�k��p�Ͱng,�5Lo>��x���ShS����;�D�l%�؉g�)o"��*횳G;��_cM٦qJ��mp;�	A����}KLO�m/�����3�*79�
�jN�q�e����e���mw��	 ��ef϶����p�׬wd-��C�����Nl<�Ȥ[����� �"N��	.G�pt��%şf���)H��ĸ�"7W`Q -�C.vH����q@]�x�jd�!��� s��9Z��F�پ�Q;Q�W�Q�̋���3h�5XcY�`ڝ�MA���Dc��dl�^���*����"�A;���iFT�G����N�]Y��)�Q9,�4�����4>�y��g�on�vN\��C2sN���"��$����������J�j&Hm+7�L(I\)_t�}(Ğ�Xf��T��j�UW�o�9��S������GGY��r�ŝK�5c+G���'-�J��J^���}�J�i��Li��!K6.�����T@Hb�#�K-�)�~68(s����6B�F˼�UJ.s�V��[�Y�B�N9Yd|���<��Ȭ�#F��{���qv ����"�dGs�0���>���i	'.xo75���aA�ؠ������v{�岽I���M�%7��iT�9�}�snX�h�7(���ѵꝦ�	ӿ��{$cŔˋ���r�����I�U!�mc�
�G��A,�?zR�/_����@�#z�^e�."�n��i:LG�����A�a�����\�{+'���?��nZo��VI��9Y,B7���@EG���v@P?"��Ŵz`��J#�T@��~-WįE�H�9����F�m��Z�R�����J7^����;"r��A���.R�@	�C�1ж����mm�\X�g΁��,q���-»\��/M�
�F�����9i���$���x��ML�(<�k�dC[n^6�Y�~���t���9CT�T��:�V6҆&(mdt� ���m���!�G���4�%8�� ��̓�?�V/+6����Z	�o����w;�[;ItݖB��aPQV�-AI���� �����n5�s>�^9��.��5��@+�,�L���Ifo�b�j��ˌ���+�����OI��;Vbb�]�q����K:&S��Ϲ;0u��3��-d%}��E���� � ʶ�yq�'#)�f4���  ��θ���,�����֋�P'��Q�v���"��KpqB#e���14T����̴��#�5��*�Pv�����i��a�a� ��gb�
�\��S�o�1���� ���w���m�iv�Y$K��&-�;b�</��fВ�R�d�p���o�o�b��E�>r��4PY�L�#�g����S�z�?{X8^��B�[�Q4��TZ    �֕�7�������G9!(�(���ZP��G�a�+^����r੿6�9�O��V���n�
��K����dBU>*���s���9Y|��!�)|4�AbΒ�1���j����w1�7��r�-pO,��7�+���ȣ��[	@��'o����fB�ŕ��x�I,��� �u�nA����DS�`%P�
9���x��d��ø*s��.���V���YɃ�)�E���{�E�JY���*�||'��N��R����"�;��YG�l<�Rt��mHS9g�^�,�a��b`���=\���ѯ�tB�w�O��Khh��~L��uy���� �,ʉ�JYq��
�y��m_�~��v�]OĎ��������� h���娼�ҁ��J�6�
�(��&����`*��<ˏ���LJ�-���{8�h����i�T��M�9�F/����Ncz�k&�b� 1I����y ki,-�p������x��L�@_xT�<���>�pM#rif��m�,�lǂ�����~���:.�YϺ#�� ���]kF𣰐�**��Q�Z��vʼ���u�D����^��n�����b�y�d���M�l�Ҩ^-�w�e�(�x~���pg���Y�G�8[3_���]��`���Nօ�>L��Hgݮ�p��Ąہ-����әRͮ��T�p� 2�:��P�Q�/3���~T�߰��^E#����<��@h�dQ�ו����	|uhzx��<��r�w?K���'O�Δ;w���~��!G�����uU0���?m,���(,?Q[
dܷ���qӖ nTt�<?�$о?V���(��P]9{}ܬ������נ���N�.�\Ov���Ǿs3\��ڸ�~ �iA�1�G����X�I��&��A�m�ϡ��-��Lq%�i�+��3e=NFI�*V�Y�7�O<9"�ac���1�L�)w�M^&�.eX �Дկ����j�����DD�SO`D5������%`��Q�j�I?����`�$��`�� �n�wet�����(��K[7<���n_11��!�%}��b3�PGqӏM�[h?�ɐU�[����b�15^\�u0J�U�V�����}�yA���	�K
Uj�>W�;K� U�܆�-�'�x%@׉HOײ�U�8��jm�8�[gLdt�h9='!���]!�P��]U6��H��j�f+�JLǛV���U��8�:�1�M�4%t��%t-<�;m�t��h*�|��=(�K�'���i*Aǌ�8�EF�;��� �8܀%�&�Wr�L~~�V!��R�B%2Q/r��dnC�k@�U�RwWב�󍍘`�sT����Q�o��,�����\��w�,&Q��Ѷ��Ƹ��&6B91����P���<t�y^���uT'����0���4��p��i���`Z̔9 \V��9Pԯ���6޴T�<ݖ'l��$��d��2��RS.��E�1��)B�7�#캊�7/`]~ ;A�Y� v	��Dpo�����*Ɔ�8g�����M��n?r?��,A}!MTaM�h�MEN5E�*��<���hV���.���婤�蓒
��?�+��1m���N���h|*W�Vjl��ԝ��;�@�/$D�F��%��=��)�I[PR��!!��66�>��;�MB����o�Pw�4>^�ML�ء`E�����v��ˑ���x�n��Z��8��혤Z����m7�=_��p�׻��{��iۣS&��%0����Z��c��){�-:��D�@�a��^��	]!���3-�6!xO#��7�.8O�Wn�eVH��j+	A%e�~� �b;Y�J�
��a!
�GǕR�������#L�y��q�`���N�~�')�� <+����_7sd��Ɍ8��� ����Ӧ%� �復�zV`qf?n�M9&H��j\H�B��MUC�5bl���eծSS�v�UӃ�^�-��nωUx��k�N���^6�UT�T���u�
h��x��ǃ��.�>$�yV� �0�_�ʷ��̧}�4O���D9Q�va�>Ww>:Pр6���O�n#�hq�Q�>�׊��jV�@آQ�Ɂ6ѫ��b�����'(rNǯ����]:AP�Ol�ٚ��h��!Ѫ��:L�P.S�I:�O-Nt��-a#5��!��M@�N;#-��=��P�O���#�ӌ
_�ĸ���#�O�n�X���;GXnj55��8����~��U���^?w����B��w��	�л�� ����Q�Z�'n{ykG"�f�k��Ō]�R����vp<̂�=��=ᆛX��/�X~�L7Y�}e�c��ƈ"��
v�5K��ը*�q:ݒ_H5/�h�(�98,�����
`�ffIHjoy"E��<=O��s{�R��H���vff.\�����ꏖ��_�^���a���0\Z�R�7�"p��Ӄ��y��-���I&T���<}@Vs����n�[��c�C@�h���Dv�=q?[q@���PVn�p�,�V=�'x����x�۠������9���V�����9�'�Ϲ���Cm�ﾜ0gq !���[��kk?D��(@�·V�D���������_r;���%�"	�I�D�ftT푪��kh���5V���-�vz��R[ʏf�29 ���G�P-�=�'g�&������2�Dk�O62V�$o��3d��O���4�߮�h5��U��dz�;Ob��g�
0�F&�Gp�	�r��Be��"���m�
�67'���':�-��;�?�D;������5XOԶ=��Y�F�^�tE���������À����h����7�٠Ɏ���Ɇz����2�(m17����C�n���[.w&1�k�f�Mh�.X�f���1ݿ��eh�Ȇ1�jn{o�e_�Pff�����6*BK'y=�97�%pO��HV?�m���A�����S�bo��{��Y=���aݝ�"V�������E�EdJJ���JS'w�_{\�?�S��K�c@�YO�RG����N�"���2�+��%���������nO��*��0�Q8n#ë����}d����@��N�TI���߀՛�&]�d#�@�9:E\�J<�k��P�r���SV)l?�t�J�����i�`#��^g窜�d���s,1gϸ�����wn��(�Q	֑-�tq��B���`ny;	�����G�kif#�A�������|�v��Y<qόi��hW�d�����n9�����T�ҥ�����c?Rz�VJ��C��:�Z:*�8�>p�h������������:Z����Y�9/y�qt}N��#)\�I���sA��+C���M�/��1�8��ݜ:����8� ���KCh{��.	��mN�ڿ�ԓȫ�r �JK:R�g�&�E�J����jg��	����n��|<;�V�M�j��ng���@_H�huc�)�Ӷ�\���OZJL-{g'$ViS�u��s��[���(qH�~��a/�BQ�$a�m�2���?�T��4��~j�B*�N�w�� ��|��OB44�TW�W���FrwӀ�z�`��=�G���vT��{�m��X�Y�v ��������E���0��1�`\����ЕA�ٿ���Y�sw���ym���I;x�c9�&�(���z8�g�_��=�2��o�
mJ���P��/c�o�gM���?��������[j��ں�J�S��i�aRTp��$��(�d�U}�ͱ�i�M�٪$H� :M/��9YO��MOM!EV+��>W4э�늛:;)�.����^�����#��z�2�����i��}�����F՞f�2�6<|�I�FJ�E0D�]q]����o��Y/ʁ�EU�6�"GZ�F:�C�e���_����ڭ���2�+b0/��t@���E��'JF~�����(�>��5���a�Ձ����ۀ��r�!C�w�����Do>���B�Ѿ�v�T�S�]荷K���$��D{B��x��UGG�rSu=ozb��������3?��*�9qvؗ�Ϭ�� �`h-o����Y@����d�
w5�B#�;���PPgS�ө7��?�r�r{d�[��,��Yq�����9k�C_�#8�3
�裣���Y8\u�p�9B\��{���}SS�B��(S+��ՄAդ�Rn^�\^Q!`�����y�%`o��Ȁ��H��<_��z�j�!����R�� ��8EޫJK�}���{��v{�_������H�F-����l���5,`nn�d�G�/iU�_YS��f�n|	�G��rҿ�^T�'�z��4��U��L-rh/���R��ɉۣ5�5�9!@2�w9 �c�e�Σ[�b&ȹ����˝��3�s/��#��?f��������r���j��y�HL귒E�[0����e���K����e,T{F��H����Clz:�Y:�'}A�L��\���ѷ�>t�P'�������xyaGiE0=��97 �z>R��{�V����1v[��CDŅY�j�$��Y��q�`���2྘����	�k��@G�ch�ur��0a=P���%�a���o��<�r���60�uKb""��g2"������|ǃ���\�DK��N���7�@IU�1��A�r�w��E}Q����C�:�_��n{�v`��kJµv:O[3wmD1���u��F���s��d��g�?��t�]���$i�z��*0 A�<f��_u�Iw��+M*���3��*�KF}�ſK;�Gr:���h:'A祬�lH?/;�.W�.����c�nC��C����K#&�e�`e�2x�᭭$�����^����G� ��j�9�}D�,�M����P�"���"9@�T�O�Z�r2g	�����BET��ɮ����9�A����
��R֨��rҧ���-��o�im}IB�ݷa����S�d|N�U�d��F}�J���
��g��qڬ&��3= u� ���d�0Q[+��W!��2Ն����F����0eӂOrkf�ڱM����7*���xLi?$d�g8+���,��+���-��Q6�ͺ-�����I�ˏ݄ޗ��v�V�	.o������ݐ"`,Ks�$���Vƍc�` �́�c6Z��TbteU����5�޴��c���N�m۫<xv�qa	q�g�1܅���������2�uع0t�d��{9d��FI�p���t��0��u}7j�nS�<�M��������7�R�T���b7��ka�ग��ww�rV^Q�`�:�N�Œ܏�Ry��n:�y�+����FDཱྀ����x��R;��b�۵��e���ߢD%գ�;~~���0c��5,�f>�����I��p�����̇�`u:TN�BB�����P*͌���5��������mZ�8��V�d8�aC_s��`z�������eIvܰ���R�qF�Js���j�VHJ�+��jಉ{�5.΅��g�/T�0��H9��.����;��<�����04+"�T�l�+H���t��1�(E��t� M�
H����A��������K�<1yvޙ{��;3��)�C�%��<E�e#'�8���8aR�%��p�&��rF+:n ��u2�תk��z�<Y8G�zEEm׉�;1��(�9)��i���X����G���=E"�\��]�UK�'�l��.޴�7(��9�88XCB"��k�s�K��Y�i���<*Y.m��C�� �x"y0}���Z����Pob�{K��{J
���p���#t9�@b5g�Ͳ��7$��%��r�~���<�II1,�8 "F�#��ĭ�<O�hm�w����\Ά2쭞��sl	���A /�.����S-Ʊ�yĚp��o���x�F��FZ>�e#�(�N���D��@A�2^��%6�oLbk��W15�]@76��)�����ߛ`�}�8I�{waJEzv�KM\X��y8�PSC�|�����������"��{�ap�M!Rh{}��cK�*zyܯ`��`�6l�=��h����V���O��4T�KW��S[Uz�}0���Z�Ͷ��F��\����g���Ȉ��9O�S�V;���BMήG�Y͗
�b\�����B�l��)���.e���	�d�~0���W�+����?�c�]��f�>4�u".��l��/����D��Esө�c��BY{|�n� ~I���V��N�nQY��6M&&�����C�~��8��i��Z���Ы36�t7�tnY@5����m
<���F_4�w\�捖t zN� ԕ%���{x�ۦF������Fb�M�� �<�=�%v�KRH�v����$K0��P����|5: ����	�"Jn�}�ίB�Vo�%�D�FF4�͓&;��c��b�a���v�${�$�X�g��E$���� �Vz�������_�NQ�����ݜ�W&����eNY���Ձ��ӺD�C��($c(A���e���3*��Rw��W��;!��b��2-ҷa�4{�xX%�$����Z�Dj�f~����V���䎼�~��|�R�����+x꠼�J���%��CM��~|۲�5O���๞�����ɹ�8�7�w�V�6�9ρP��уM���cK*@b�\�޶i�FX���������e!h��G��g �а���΋�~����\�t�wYF?2]�n �Cw�� ������Nܡ�BAT��è��1i��k?��B�4�`[��W�S�VX��ş?�DϽ2޽��w�����%��|,2j���w�7A�4���S�.���i0q@�忴��ʋ3����n�������U~�y��rR�?�u�<��tK86�\́�� �ŠF�qG�/�q���Iڻ�Ѫ������b�pY
�i���,MH�����X�Ngv�::8�Ļ>�h#Z�c(`Svt�ԥ��͗rv �Y9����1�-:6�+�Ӝ�֢�Uz?����0ޟ��Y2�K/�;.�=&�.JJ�Q+�#���r��hW�:*\ĉP���nu|R��=��=�cc���o�'�J�?w!{o��H�YG`U���R����镏?�����;̨���g���z�6B�6t�3$��A��H���zA3 �9O�C�.��ď�њ����ƭ�p���}�^�w�ѣ��	7���~�Ue��BM�:�7q�8�M_P�C�(���z��_1�� �˾�����'G'wCf3ʤ�F:Kڒ�E�![�����әz����W��Jf�أl4ZAbS�4m��)�[����/~{m�,t1԰��DD,��� U��7lGߊI�Ӳ��~�	$�ݸ�b����B�L�q���É�)�$W<}�i�����	�������"�b�g,��Jk˝�A�"�BBaP���q��~�x�4ָl�������Uh��SK�N+�<�m�r�P:,���J��ԫ������O�o��DD�c��Z�g)ҍ�I��޾�I��g�n�l��r{zvFYY#D4��l�ф�k�%cÊ�S�XB���%�n��DKn/�I_9
�+Nc�i��79�v}�bB�ϲ�l��m��`x;hy����T(��~�$�c1��Wc���S<W7;&�s΁Mk�Ub�L}7NL0�	��(}\nQЅ=�LK�$ߌ����c���,�\Jܖꇬҿ/�EF}�q9���i[93[�~�mj:�{PԱ�d'7v�
O��1}�TDa���HQ��F3xz�kwg�����&�R5y���$%Y��D��(����R���y�E���뫿�.�hu���Yƈh���c4����Z�����߅�� Q�,�8�hП��� ,r�5~{�:!�-�����}�+��K﷋����GY��E�{�,�P�r�Z�µv�ŋ��ب�^|k�����!���{B�r�7~��a6 �}u��Wbj���2'��vᑟ���i#����ST�X�"b���~Sîo�tC��X�������jf}�lM��a�E_p4Ɇ���y��Ҵ?�N(Ei��U��B_Q�Oo��5�.0?��W236P9�C>�x���.�_�ca�Eu�67�i����Q�xz슼:�|�v�7�_��
�Ѷ�[�|��xVԞ;��^H�w���C���Ӿ6e1[m�0�g�s�P���M��4�1���`���ˁ{��l�ҋ	� �� vP^��	��aߠA��K��}���8�8�Gܹ$�^rcB��2�N�� f�u���%h>���EW�a�i׋4p����Y�G��^�Ǯf-�T��������}y=�,�*eVQҟ`ө���q�$���q�w����@�����Bm�
�l]����d�%n����s�COA�����8Q����x�=<�u�����\'��.�	�JI���z�$�t4�5Q�_p��!�=K�|���W=v�K�±� ��cg!�]�~��AA�����B���6�y�V���w8(�Z(��V6�额v��ފϵK���K�Y�|�1Rػ��ߎP��r��&��P��<����갈E��[�t�wD����I�;�jF���yc/Q��`+K+2�h��\
��.���r�:�`��Zb�X���ŚTib��xgB
`�v[VA+t����]������@��$*��ǆ� ��#��.��.��準}�M�!hEޒL�3"q[�v���e�G?�D��on4A��V2�(�qlY�c�(��H�L�,��]\�֬���i��¤z������4ɫ5T�&��wYD���:�z��O�W�l��>�P���W���w�S�I�NPV�����p�)tDu%+��!�}�F���l����9����:�C_�p���Z����z.��n�J+c��ӈ����K���y�h��
�'6�}g����@f��������=9�K�Iv'�$L��e������]�s��SB�y��v�E\�7�B��wJ�}b���E$�4"i鸳�O�r�������Ob�:P�����B��v:��K�	��@��7�=>�m(�&�a���6@E�r�E�c`��U��������E�ӯ��h�B�ÍEZIc��RwG�s�S�En���$]�tjrD�n��Ŷ����=cά U_tɌ���&@�b88  q���Y�F08���1�[ �x|����x�;�-qb���'���us�Sn����q܉u�n�!dkϰq�~��e@�hlh���Ǣ_�l�!:�㝇�����K�8%o�x
@�����}~nl�!��L���'
���5x�����|a{SY��2��gP���x	vdа�	w��#�IJ������ P�`	�-ЗM�|�����	�|�އ�a�e���u����c/V�b�ޙ)v=X����s�oEm�6���H��]���aUA�	��l@V�h��o�$�l�/���^_�����b�+�;��aE�oT�B��zI�<7N��йW���.��Ad��V�i���ǋ�	2mHY3��g�+Z������
�3�,�;��I�d��N�L�b��j{��
�y�ڤ�^w""6b�������;=�e짤Y����*gAڙ/���9��J�d�
�ׇ��7{b�ݺ��,m�1�Qo�8��3$��g}5?�H���WRc�G�ñ�i�{�(�-�[��������o�h�q�����[F)��H�[����|�p�������E]�^f8���+t���M���,9�H�[�0���twgĝH��-F�j{"�w��B������1��� '��I�c��(��;eq\��zn슈�d߾�~�;߃?�z�J�=I�'�I�[u����F�XП�9��\Bͩ���g�T�ywR:���\t�K|}����j�7���[i_�/ǿ9_^��~��(U�߳�,ӉKK�Gq0���b]�~�u����:��k�]9#��P��Y�������W��}T��y�:)K�rDq����܊�I�pɩ)C��/�6�N��a����5��m���}�����(K��ݑ1H�1�����1���(Ov��f�!{��N'zZZ�o�^��l��N~�f�:�%�V���B��VL�J.瞇Ǜ��vvq�g*��abd�	"�����������/0)c�����Nn� �8��muu���J��׆�U��h}��W~׍�.;�z)���\����\�f^��4�;{C����;�X�C��xx��g���k�՚[+��{�k�n�̺!V6�T`��n�f����;�\��.��Ǝ9��^֙�n�*��h���k�:��Yп`=g�Mu?��I2�d9,'�z���/���3H�����#�Ǚ��E%( 
�ru�s�%6v4OsZ�/g���۳5��s+���[�Lj�}�kS,��dh?���&Ox��;�I�����ۛ����[[z����AR&t�_ъ7ܰ�H����/�t��%f��l����Y �/`E��9�}�DO����
�s�4�W��g"+���;�j��>p��
6���ٕ()��~��m��{E̋��y˓����V=�է�O HF>t��k7VBkC����|��lt$: �����⢞5=�^o��3��s�Sw����hh�Q��`D�~����C%R�O�I��SzI����/�wϊ�UQ=�?��c'+�$1�U]=����,��ie��L�E�E6g�To���4�ܲN+��%g���f�x���jT��-!��ِ�	a��C@b�m]~��4d���؝���[�f�㑕�X����>���a�m�S�Z�f惆��U�"8/8��s�	m�<���j�}���W/��m*z�.���{t��H�-A%;vT>��JxR2��;`�귳	ņ�ev�~�	�q~_���oB����Q�3�x��c���'���*]���#��s��I=��e��\�H��z�t�D�{`��qq5!���ƛ��[[�7���}1�ЦT_qZ�d�![ ���!:�F:�M=
�r�D���ya��{����b>p֤dۑl��#�
�K.����=f��*˗"l��j��LG�:Q(�V4��^i�S��s���j�
 <��rH|�r�y�
S��9�)G7��[I�81.���\�r���'��tXa�23��c���dLA��s ��@����_������X��P��CF������b�B��)�az�J"���ޮ]#�{�����)�Jzazz�;ү���1����e6zU���b����i�&��ГD ��I���,	�.$�=�-���tR��q��{=qU,H?|�1buu��S#�T�;����R1L���g���]�Nv �Z��]���;3P�.]:�>1��nn��Y�Ei�fxlF�������glc���:2`����hii9mp����?.FŒ�O�f�LHg�L���Q��<�J@��T�\���V�(��q��������8�
Б'n-��e�@��<�ttTQ<�~un�� ��\��f�O��.;�0 �^��YR��[/����BE��@>(�����!?�ʙ�X���`2p���LN]��-��R��d{JiΥ%�j�T�eS��[Kg��<�cI����gYE�ͱ�Gy	J�(���c�r������g�q�P6X�)�֎���W�e�o��2���'���
�h!�t{ʷ[�����ji)�|��D_p��2RZQ�ޖ����K�����1��s�Ʊ�_<Y0^;�B��rF�Ui<�.h9ʶvׁ�O �z[��H�ue�������@!Ʊ
��������t�����LT���U(,�b�l�uZ� Ӳ��'��S��D���e�Y�by=T�ʆ}M��7L�P���^�D�d7y�CK�7�-tL�s������*�p'������;�&�=�_p���%&g�z�]��HG�Ի�"��O=����E7<�쌉 R8�<�xWZ�;�S1��Y6;o�L/���^���+�4<�|O��ʟ����-��N� �(9ߖp�0S��vH����5�z�`e&������_j��E]��s�<���/�Ѽ���o�<9!I;���k�n�$��	~��J�5�os����'��Yz����O(p����J)�BN��+����iy��4�O��x��OcO�r�lU��'��3)��f��q,O+_z��������Df�{��ŋ���s����\�k����]&gr� ���u�8\y�I��۝�/�
���lw-31��c^���Y�l�kg��L�D5p}@*����'�C�>*�;��;���n���x$z�d�\��ރ�F����迟�p!�w���n3��N�jN�-��q;��--�X������
O@5�O�;�-�T����_�� '��?�ݳ�Z/Dd󪫫���������uV�Aa�S����[��k8�x�F_����B�}���
w��P$�ܾO�La�����KYpt_!v��`J�2V}���S`�Ì9�|�n�dkk����:wGf�ckѫr������r�>��+De�r���yr���ι���oPmz��g��Rl?������(F&8�Rן<y���]�L�P�?����)��%<�n|{>����.V#�u)3��������wc���*���0[w��H\��r�v�7�P⎟�u�x龳�qϣ��3���ll�f�F����������P3���n<<�{�>��j�৷�{��F���\q�o[�ך���0�xD�s_F���dV[�py��p�YeIx~��}L.{�c�+@�
��{�(-�]�������_�گ����U!8�=H�6�,*}��G�¤�5��72u�0��E@QY���%��d����C��Y�ɟ�VL��G����u
d�l�ɂz��FNm<���o�wv�Cf}��Q+��`J�L��I���c��
�����Uo�d/�=�i�4�?��m�;�	��$�ہ� J|�}�����5=�&Q��{�>$ܿ�K�����aݢ�~zN��rp؜i����hw��`��W	uz��&�dJ�^�	����9y0w}�,�ujj[��B�� `�U�@Co�����R?}�յޥ!lV��ى�����N@�̎+����f�N�T�k�k ��ԇ��1��^�R���
�z+�ى��Y��~Tbr�n�e�&x[`��j��!ڌ!+:2:Ҳ�>:َ�l6 �)��th^^���/�%�ZVɡ2P��[{��܌��q����FƝ�(B}�˪ߚ�D�����K6N�m�S�,m)<�Kφ޴�c��G�jl�P`����� Ս�zH�'�����\���:��%!7�^�A��5){	G�ͮ:g54�DI�F�i��䮍�,�s����5\�����>4] ��5^%S��̂9�k�\�/�~~��R\PbmTI4FA'm�`-t��3���˛��V�_��Y�_v��*��d?On��b
p�����f�ڙ,�yъߏ��u΋�0~ZIួ�_��"�W��ɧ�Ɇ��%�����p�&��p)�N�k�\T� ��L�Y�O�h�k�0����`����:��:����$���jݳ1�N�X��~���Ώ��q���S���hu��)�)j�hE(�XF\xc�g��d����I���TUB�o^�d֎��γ���&�4��tB�����q��=�4�D���q��;&�AfL���]a�&���׌�ǥ�����c�y��b��/������'�>Ѥ��kA��T.��a��m���mk�D��޲�#7���6d"�=Y�����I��|H��)�U?��\]���@T~�诞�2l��	>	�7Hє7�>��<
��R2�ܵ{�>���#4��~�`<��eq��+ O�U�����z.�����K�f^5�8�#���0U��}�Hř�h����l����X�M�9)�Qm��;�B@X�2�� �(���ut��O�n�X�SVey�I��x�X����'+�޸�1�%��'ՏBtXW\4��B��Y��B�ж��n߿
4m���1<`����{�0�l���:�Rl������=�b-�;[���� 16��Â�.��=���'�25--l����D:z��~ �t�+{�*�R"I�3t�L ���yo�n�"WA��Lrb��Mw%ŵqS�Yk"J8T	�����TH�uqTYzل4|�V��R�ʷ���N��������;�I۳�j ���<�P��Oؤ�6�	4ɏ �`�E2w�9�M�09&�5$�f� �/�x���AcU0=�KֿD7��Y$�T�,��31fZ�z�����G��T��Y�2����ۇ�y.֘;�/%��+���V?������z��cGPt�vɪ�f���E��^Jn�%���(��0��'�R�}#�x���4��+.�Z�i*N�7����̰�� }Ķ~@�t$j8�uu��s��ot��b����j(tP�
�����v���Y(CM%������l�A<���3���I*0����Ke��~|�Ě6;eXFHX�%=��:��0^��u��|�77���:�;�w2y����R~�}�=�J����/��9�Ǆ�&�:�����熁 U�m:3-99z<�z���,��I�}�3�d��Ϳ�l�D�_Α
��>�I��{|V'=�1�cEsI!�����SLv�=�Ӝ[<<ڎvksKdU�:8x�Ib� �t#I.���v���,���F����\�q#'?l�t�F���e�܋Jl��ȑ�`��JG#4�̴�w�����չ(�F��o�d�bɊ�2�PUˏ՞5K�а�N�� ���h�}����;�d�����
c����G*D����C�ڂ�ΚD����.J��:�(�7If��ZeЈ񽖞�`�G���z���݀$/T���k5Y�h�]S.�k��׺S�A��2��BS�����&Zd{|�@mf�p�t�c�7��Β�Za�2Y]|�kG���#��[�����k�Z�BY��G�=�Y�B$����?��rK~�@�g���]�9!:?���><y"I{��{��o*��l(������9����Z��[U5��m��v����)l5��������#�D[�/{guly����T�r�!Ŕ8Ɂedu$d�֥=Uq]���;���'�����(�c �?�
*��Ř��,����`c0���g�h{����6�J7�ZX�,�Y����Z�`j����/�O�J�B	ސn��NlO�����_�G~9vz�TQi޲1�9?���J��:J�c ��Z��Zk��@����=���;8Buz�s���yk�u�=�5�����2���S�5����ǩ�3;ĸ}�>t�b�J�Q�F���.F̊ X���°� (n����{*�M:�5��G=�������}� ��9����(iQ D��"�-;mu�Cgo�RhV�ߓ�(�9�ü�D?���vNn�̱$*)��k��y�n����ٓC���I����_uP��� |c��W���f1�/�~�@�Oy�W=�tg�J�5���)��Ϻ�=9��J�0�-���	��&ܤ!
�7?'�
^������O�.���X����R��1�ɝ�Ԙ�r�p\_��Dׁ�]ļz����}�S4N ��C��3�T����iL<��Kɟ�53��+G�����}��3�A�����n�2~͍_��ؒ�	��ۓU>e�������t2 ��Ƶ-�9YGM�VV�\e��
I�~e�>�2�g��������tKg�f�R��=��w9������^'��_ʌc&�����pL����<p�A򏧕2hF᡾ӳ?hg�=�����P��F�������|�:��<)JT��QT:�Qgu���ֈd�հ'�O����9N am� ;]�����y]��l��&i�t��px�t���a����
5E����OW��q9�H
<�k��5+h��>�{4�o/��Q�2rR���H-��2��!�;S�
~��f��d�7���ﲲ�j�n�g�
�~�V��+@k�A�駲uX<��gB���c��y�¸ǻ�y��C˴����Đ<0w.��Z8E[o{����[eC����	�<FX��"��3�?��H���_t��/����5 ��ޢ_[V��7N9m��z��Q@� ˬ����� ]�M�����vT���{�RmD�ZZ���hG�9�b0nyp��&I���x-�$�R��{��;��?����7@M�{ɟ�#�i��"g�2Z���5�f��\�d�\��1�pNR���7��'�s)�$�<�5}���ĸ6M��:Ĳ���Ѭ?K��>�$�o�IZ�\��E.B�jw�~�2�w�A�s^��z>T�8�s�.4�RH�S)�f�s��1Vso�`��]�����Zo��[ u����"�b�Ny�M��xΜt(�����P.���
/���T�&,��T�&&Q�O��(�};��fW���NR8�*��~�U��T5�h�p�$Q:۞&�3��c�݊�\A�<#�\��ҋ�}Sܯu5y�m�~�O���I���X�������m��]fΤRCw\[�I��br޵�z�Rr�����L^�*��׍@���iF���^��A����;��r��E�XO	����)S�+��D�,�����f��=R��A�`Y�u��ʊ�cIa���Y>����V.�XTt�Uu4�@m���)�Άh�*���$���t�a��[ź���I7b�|��am745�\!��0�!1*�f؇M� M�1Ԅ(�e.��"p������̢$�n��t�.)��Ϲ������OZ����� 9����SU--m�,��6�j�2�'�������E6{�<bWR��$TB����3c�!���mf�|^-ࣤ�{�yN�8���P��ռ\��ڛl�4�Ɲ�P��c��#�r����#��t�/�u�X5u�8���_0�9��x�tB�)���$��<My�tzbׁm��z��1\��o��y=�/�7͠Hr�������mr�2��c^x��˄.����ܪ[r�:�jYd��
�=�Kj/\��4�|���/5h��Y#���$�� �aZ	"�S�f����a�kT�����ȣ�W�ːj����&��� �נ�4�v�u�_�O
�q�7^ⱆ
�����ퟝ�j�մo�BCE]qmZb����_��0���t���R��-�n��P��Xz�VE�_3{�Bﰊ���/+�kn���-K;
|D_��X?V����6w]��2d+I�t��9��YG�t0y�U1)�W�Z�LcW�l�+�a*d&=�����$�%�������Ը�C�~�T-�+� j-]�L�e���G�/�9e�~��B{���1��3��,��?U���"��@Uq��>ˉ�����V!��~�#x�\��(bk�Y��W;R�xdU7��7�w�7�����CЈ�a���o�1)�܄̺�h֑4�Ƿ�"��)�v����2U�� q��^�~�Z���8tih��
{g��0�����яJ~�&R�3�&��Y�PZ]�/[+x��i��&i
�U�Z��:N�X2��.^����5���,�T7T����&�Oׂ�´lf:�I�f���N%�8�b�@�}�\ŗ3�]�ת������Y\Uf�1�b�k�A2IU����u��K��@�n�Hڱ��)Y㏎�M_��B��"����z�Y;���;�9J$#��%����7�W���V>5=a�@��뮉I��Q�ba?���[����z�x=��{��
p�R�X�p<�=-`W���+�f��k%�ը��8����`& 7�K|6/�a�u��u&���{h�Q�A�C��O)rV�9{���g�5	�]�B����<������z��I�Kܕg ����|�O4~U���Q��9�����*%5U����Q��JD�}�M�ζ~�E�0YB�2�0�Y�"����U3�_��0wD��.���H<��C�7n����r޼�����]����[���b#;��8~ Ϗ���G	ʧ���x^��l�Y�t
P��vZ0R�I��u0P�3�q�I��+P��Е鳓��;e4�R�|��7�)y�n��)Bmi+�b�p�����M��+��b�hS��(E?�W�@�2H�3�f��69d�x��T�m)quw��=rcW(8f��=	��saw�9��!v�ӕ�>���U#!�p��t��t�\�;�H�A���?� �Oյ�~с������ /:V ���!��	�� �M�� ��/:�K����er�	q�o��<��k����ʕ�m�1-�M�;�0��X��)����c�S�$��NO��c�V����,�8^���;TYc`���?I�l%)QJ86J�id��킧��%�'	/	��ǭ�t�˟9�L�p�F�B_�G��lx\��\�ЬC#��$���m'��vr��g�2�؏Lk�i8�a�3D�;;J���AH���p}�d���ܢ!tx����!F�Sv�/�q	I���8B�Q��K�����1��ܾ3����79HИ�[׿(�IQ�a_Ӡ�(��*��B3e��_	gg$a�@ө��4ŕa76nȏ-֙A(\_�2Fǂ�W��?><�ڎ%|-H���4e`�)���������E(��zw�ʿ �ϣ������t:�X~O�zl����|��K�	y� ��ǎj���}�f�Ȫ��9����Wt��xx�z�>�����>	�c�Й��P�4ZH�D��$S�Ӕ�v�L�+��T� �l�; CHe�26f������jH�(�=X�b��~i	I�A5�g}^*��~��i2�De+���Z�:#�g�Z�v| ��w�*���mm�>��]U��
F�D��ȩFG�c�r.���L�v�H�Y��Ҵ�n�$A˅qy"o�5o$k���K�B�m��<}l7��+.����O1�Y����\W���d�ڕH9N?m����]Ԣ��o��� � 6���E�¢��S����9$��=+Fɟ�G����;?���ݱ�OZ@�ˤ��5E�����B����]+v�r��;s���=�37��!\zj�q�!V��Z���� QAxw�{�fv��k�<h�C*hXh_����~��ס'�w�J��ì�Wd[�?�� 1=(�7�g[dϢ�6�p�j�|���ܵM�#��抭�f��e��JKt�,�j������ ㎉�R������PݐFu<(	%����҉��!!���`^��^+_b��/ժ!c���Q8�٭�Ns��P`����X����?��HR�+~��(�����s���ruU�`F�q���of�D訰�hJ�i��'iә� vzVA�돾�e�ȡ[i��n.Ls�GZ�_�u.�eQ�}H�Y������#����~�bͦ{B�!$v���u���<���m��kSe����{hv{����M6'4&F
��_�]�bg.}(AR�����2V�g�Ũ��ۨ���T����4yQ�=��yE~&�[OOl���'._����'輒U���G�k�bI�	����ֿ]�7�Q�F�D��8_�+~hS��>j�n__�_B�x*���X��{��|��
W�G+բ1��䕭$pQ>=,漨m
0���6_e%cbsP�t�ix��	���Z�c.dޢVk�p�t;�����(�#*��Bw�f��+I��8� "-���L?J�O%n1;���O.e�㭓E�}kr3�	Ð养Z�E�]۵�E��!��u�Yl���*/pvd�|�����Uҡà���*S<�Be�Xۓ�@�+�zz\��?�6W�(NB������|�f~Dgd�6��9�-�Ф֬���2�b�;��tĹEl��O,���NI�8ZLH@��w��f�H�4��j(f	(pY,����
��e��b�U���>5��?
�a���o�jYK8:ݕa?�l����l;q���z��G<
8�<�JH����,��!�z��&��nvV/rX��r�i�(�.n��N��RT�^N^J7Q� q�����X����y�c��v�,�T�^rN�F3�J��j!��9(��Kk�k����,,(�G����׫��	��.Z��D���(pPp�(yܛ����h��:5v�;%����\�[J�Y�z��͞��F��>���K�e�+b[z�U��L�������[ぞ[+�78�	Xg
%��p޷i8O��UX'���_
$�+����ιbpS�e@�-v�y�Hq�>���tK/ը�-M�Rl)_��w�D��G���3���� �*DC�dX�i�5�}
�ߑ��ӻv���@�������d"I���x��p,-e+�}�%7�%��t���@�M��3B:����/�2��&[�M�����ݥ�k��H��<��b`��?�3����4ڝ�S�6��/���[�w�2Sr��������i�������oƋ���l����~�M�S�Qɗ�.��$���n�*����M �c��ڳj�2��R*�)3�~�+������yQ�_�з���H`�	���C���_pS�znSƘ����ף Ni��~ee�)>��5�����Lp7~�\S݅ϑ��	�c==2�(4�  ��e!q�UK]����BX��C���#�2q�τ6�1��ץ�y������eFr'��eĔQ.#�d�LtR:�!�t��jj���֯�F�ʻ�����&T�v�K�-A��C�Ƽ@]��V�-u����`3�c�އ}W�J���C|�3e`2��Tw��T�O�����-�>��,򔌝Q�IT���.�[�Y�^�4�=��@$��ɼsk�EV%LɎ�4f4E#�/"�;�왻��T��,���L���>h�H��";�"ՓX�-B�d5��Bůl{�SR���^��h�� |\�?�u�Dȶ�L<Լ��
�%6#�h��he�*��0�VA�DMK�Rh��?1�I~�c�d��a+� ����3�C���m���5]ro�ی����F6�ہ�7��J*7��մ�A�y+��Kd�;�UV��:[���Cv����[-���l��6Y���q@kq�;.�ٿm~�C��V2�TL{&�(�5�i_�CH�Q�`�znx����o}}���'�� ����R������q���Ld������:��r�Q0��L�(�á�#Z�T8�Ax��Z�fߴ���
�d��]��� ����~.>]A����-��7əx�?��8^K�C�	�^d?����ٓ�1Ɵ�>On��2]Wa�t7�v��XC7�%����m�p�Y������K
��B+[S�Xhp^T��v==j	,G5��K���Ȼ�7���)K��� <����;i��R�f��׃`�׵����BipK5���J��"�UW�xee�
�K��L��J�m��'7^C.��V6�������rAzo՗���3W�[����kP�p�-� �/ϧ���|�uE�!M\7���x��8��y?C�G�����7�"W�֢(R�@[�����s�Tt��O�3�o-�v�.����?���c��W��ixz	�j������ŖD�0�V��n���R���<��G��O+�8�>��?J�F�a}ZV���b3Y�g�e�uA��������.��@��X�_0x�������8�tZu���L`;o�f[���_�Z������7�s��lf�m�s
��u�ض�"�"�DF؊���z�kK������dy��0E��(������3NE���F-\�����!��@�K�u�C�k5�%cL8I�w��W[��:}��֕�]�>_�����&��o5S�j��\ƞ��}���*L�X�,���&����W�FFg/�≛��+ywH�v��)����syĖ}����x(�1`��c���m&
�E��5�<�6xgL�����8�'�2�7��kC�C��:�R�u�_C0�{$=��Y�3��T�`�9P��ĀGd���h�'�a�D(3J�.g���q�^rn�}l:��Аʽ[���%Z�#%*�!�~Ҋd_��b�?xT�y�-|���N��J����+e����f�c�#�(�tP>:�_+u�~U� �ԫJ+z7���<r�:�1��v<���1m�.x���'�	z�{@�������)q�ʘq�B<��M��J�H1��O9�"�i�=���^�L`��9��������_�	F�>'?����L�W�KЯR��T�w�ק3�KL����=��ոI���q7D/�߻�~�Oi*p7L{jJ��0�pTU�OMk��`�p�_��������C��H��@V���rm�08s���!��WP��-%HR\A_����h#�6��Y�UR�����#�+e���C_����bu��@��c��[(K���GШ��M-,w��7���G��z�o�N���N��(x�:�}$@�,�%��B��
�V��0n��uBG�#h����\��݈�����zV�z�Ks-�<�QGEr���Y����_�b����(����{�Z	���G�@�263�22]�1�R������d�Q����732N8����yq����E�<Y��SY�B9]Q�6�ua�(�!d+�n��c�W���~jr&8�T�y\���E5o6��0��D��nd��4�5���'@�D���Jp �|[��C媟΢4�8��fYV�H�z� ����X�~�Y���!���G�mO��Sx�U:Da���3�s^���U�a��i�qq�Τ��r��jL�Ī�$܎hT�v�J�g�pJ��J�f�ػ���I�АL�oϻ.h�d�p�r�	��5�j�u�Q��1���E�&���\��N��$W�[�E+���g�n�`�W\؟.X���c�Z7=������^��M�uJd�Bb��{��G[R�9Uڌ�a�����g�����S[b9V�=�$��#Ѧ���CѸۋ�w����T����_��gD80 �_NNm���VH]��q��u�E�޿�#�D����q�P"F���P�[���
ݶ���L����)Ӝ���7�n�J�@��Ѕhb+��wǒ�����A�0/���#��?��:q!�q��u9��o��yH���Z*z���'[arڎޢ���UA�s���hiI,3���/Nr�&-���V!�oM�տeR�ra������fz]���~��B�QJL���Lph��=9�P*���T���އ �ߦ���&��u��Xb#�0u@XلQn=@��kCUV�9��S��y)[������G��iS�6�9��`�a�َF�ov�g�����X��Δht /�i����W|{���ѓ��U��O�`�t�Q�@<|F!j��ڶ>�@Ql����I��O6���yN�
��V,F����b7-�6�Urlڡ��Ș�bl=����2���)�0�)�f`���B�?��)��A��Y�bܯ�W���ܜ�����/�E]�׹�Wu�Tʓl�{yr�.x�����_S�d9�q�	@������!U�lo�rriZ�d���N\��o��j�A
��Ӷ�+y�}���f��.�𤕦6��P���4mA���J���8�o15׷ߘQ{����g��+B����f�-D���TuU��J(��~G�cͪZ��/�Ñ��*�w�

ȷӽ�3#{݇��El) �ԩ��P�I��6�U8�Y��]�Ԭ��u�7O#&F��Κn��x��T��a��Lپ�
j�r3-$1�e`�O3F*\��xk��|1s�j�P����)����W�9k�U��n��)^P!��;�w5w�{�8����ܔ_��=�t�pkm�?��ub�O��^�WSYv���׺�_��l�,Y�ȩ�pK%�U��@���-�PXQޤg��Kv��v&B��b"��Db����ֿ3����ן��X+v]���R��uo����������TQѤ�o�I�Y���O���"z���\��bF�I��DǏ��B�ژ����"-�}�|rj�����uX��]�Ol�o�ҁ&(���\wj19'��M�~�ൗ����{s��'qW���Z4b8|�<J�9<���X ��E0��3>�'D�t�If=���(_��D˵�>*���$�����+)X�Dɓ>N��goN����%�M�t����Ì�i�������`#��pYb��;���D�n!sdij;V�����_u����Ct��7��2��F䳦�4z��K������Є��gXTW�><�L,hb C�ĂR�EQDA@�h 齏�"
QF@� �m�H Aa�(�0 ��9�P�������z�"ל}vY�^���>� �n"���'�U@�ʾZ:v�%?��y��RP��O�WP��֎8`8<����5/�Η�㖜��'�_�a:ߕ��x4��"ںOf����{t�ݬ���o8�_=%�m��a���{�R)�ڑ�F���g�:T��(���b&������M��~]/��HO)? �-eB�C�W_���*������9t��S`���s23q=#�r��������E����M�:�W���d�<_�5��Dj�n[
�����X{&���c{�������%��,�oη�ǁ��Q�&�������;I���I�\H�w���|-@J�I�^�e~�Ț���F�5_}mi-6�'�o5Rג9��ۈ��Gm<�J�����d��x���,�Ǔ�!���ڗ{L7�ن��ʸ����?Z���&�����?���촡-_�<K�(_D��DSO�.��#,�:��]�'X�]����r%��ȣf���88�v��B����qX��PVN9��&������쩆I�0�}R���>���ށ���U˾E��X��E�5lv����������M%��eiE�ͫ�qgG�߁���cv��2�އ_5d�tD	l����ui���g�Ԝ�-E���j�W�*K���`�����.���S�/L[J�XK�d��o��� �6k���b��_��}5����� O��{��ek�d0�mW������=�'^�l��A��F��eo�5Aphg�Xm�0�'*�!]˞[�R�bd�>�Y�-̊z�l@��`�����}���>��,�_ԏ����gfLp�>�%�ī,�̙z�j,�ZA�/n�z 'Q�<��_c��eJl�hRIե���)�0_~x���|���=tl��ޗ�G��� ���]�7EZa��N����}�-y��:`��:[}K�} M�@�N�"��	�f~žڠ�;P���6}�}�4���/����ν�Ik�*n�+q�����=�l��� ']��_\=Gݽ%��/ᨹ8��F��kL�E1��d��:(.�w��%�l�M�� �����]Ăj��d1��fy��l�p�K��2.:�������U�����_�����w� p0o�֧��(Q� Ȧ	�����ꖼت���b��~����N$b8�nT��$�B`����y���h{�I��]��?�� �����A����3Պ�pG}�:�p���GŃ.Hm�8�� 4�F��+	w�VD������oF��׌!�.4H��3��{�|i/�S�j!V��)�I'�5P8fʔ�a�t���n�d����~.��b�X(��_۞����KY�)�P.��{�h4?�^���d��
�N���ehz%�pt?�|�'�EA�;Tc���M>��Y1���"�/�&&ZР�gao���ԋ�Hi��EL�?���DYc�;�f'4�
@ɋe�ɺ}�)�H������5�t�������������g���b���;�<� WՃ���noP<A@i�'��pbq"�jwN����"�[��ͳ�a��%���������]���/׌�����J8�p����K��F�����G9��v~^%�R���+�*;��W��N�f\��,�n�!ע* �_S8z�'��y���`=p(�b���mY����:q�*�/�����:�">}A��˷ѧ^�u��MU٧��4���?�M�iz�K<�~:��]�?E�l�,�HE�.�3�����2UZ�;�}z�X�����Gf7�K�jX����ʲk��	�3ypFx�|-������D\r[Oe���vԄC�L�u{�Ꮏ<:����^I���{(�O�m��9�yth�O>6�	j�~��Y��np�}�9p�0M|^��X.����X��	��?��(�����`4E턬���.�+O�{ ��V�VkBU�Nm��k���3��gW$h�ݶٍ�耤k#�� ��ϛE��޹����g�oVs�����065�0�9Xv#��O��	k�}��9 5W�Y�M�����.[��w���h�\r)�p]F��O�M^ �tw�A"���v�×�0#�P��D�n�m`M� Iz���T���0h�����Ur�HQp6��7�\wo�<�TB#�O��q��U6�����,��znE�_([�G�L�;����ǯ��N����paW]�G��	$ɜ"��%�;��g3~ʓ���K���eb{�p�숄��yW������(H��N�����p���D��ǧ�׽%��_���p�ǃ���|V�P�~��k6�/ݓ����?�ޖosd�5��'zڏSv�	]�s���v�����*�P��ۈw�P/����vן�_�zۉ%�`"Ur��h���x��J�݅I�K�vd��qw6	%�H��B�n���E��˚���;TE@�S�D��M{t<��I�&�V�����F��
����u�����#�J�����A�a
�	���6��N���c���k��k^�X��m#¹kǳ�XڂMBW��{_��_C>Q~/���K�g-K���� ��� �&�r	�G��������fzP)K��;D���A��a�9ɪH�q��|F����O��r��3�,a��3�"i<ǵdP�ZN���Hwp��(+_���=�����ˑ�7�oSqr���dm�+X�T�v����� �+�={5@"0?�+U��ܕ�,~�qy�
�,y����>�0�܂ů ��'�AcQ$]��ߢ>?)e��ζ���uo��,���kk@�� �Zܾ�����$R�B���/Yso��;��D�BN{������2Q4g�/������~Y<B��kO����GQ������ϧ�g߰:��?ڊN���q���ώ5��;��9�+m��yK������L�ܼ���n�r����R�D{������C'/�n�X�;����;����;����;����;����;��B�9�6�R+��л\���^���R�pE��͉K�..����쩝�L-|A�U�v�ԓ�z�E�b�'�%v��7���^�˭���{���{5�ސ�CGVZ��7l������]�#���gҶI$\{�LHw#ZY�c��YI�Q!���5x�H*��n�L����ZH������˓�2�F����H�݉yVf�n\���Cs��"+��u�_c31����1��59g��_К�o[ۚ�E��_K�NL9�ipTCz;6���s�؊U����չ�9�>7��\;�ҳ��h��Qd����T��엀�t*�0�X�Ŝ��>H��A��-g�t��-��5#��5U��ji��ġ}����ڶ��~700�Ԩ=ňgcx)����4�>�0�9����1g�,�,��Ф��ϭE�@eW��n�ų́�w�	��~^�۝�~�`O/�R��k���w�㛨ў:h�����ō���bK������:m�(�AJ��F���Z'�/���G|=N�̍���^&؍��/=7��Ԍ��^�D�@��r3�h�|��G��|�>��a/7�� \5������2�ǱnV,i�	[���p�# �m2�4�B��o!�����	��k��ԟs����;rK�ml����er�#2c%�R���̹�x����&*c�G���a�Ka(ֺ+1����u�-�D���^��v�z�ў�6[�٩��Z�}2�VIav��E�;̍�A���I��w�Qsʼ:��b��.�� �^ݵ�3e��p�թD��;i7n�X�pw�d�o$�NZ�9c�!+pv�>6
�Cvp韮�������y	�I�#��H&����VWt2_:��1����F��3�a$�Y�Q7�C��2��2!v�LW|� ��t��v�;ג���l6k�R`Ppg&d���φ[�:��������S;�xǟ���j��[v���¹�Bn�V�Z�l�dH�GG�9�82��ue�w*C�2O��p�3��qj;����qP�ZN�O3{zR����-��+�z���n�[�F_e�AO'��|.E��M�!n�K�M:Ag9S���F�?am�1�rN�α�8hNJ�_|�]bE��{�n$�������#}ֿ<�=�>�(�����ư�W� ��eN�Bz�F[�#���t{@�����,.sl�+Q�[5|#`���Vy�"�-���=���������ߧ"�=:5� ZX�$"���9�'�{۾���4J����nΗ?~�reB���pe#��0 8(�}��a��֩�وY����~��'�2ݹ�ΰ���7����C���|�餬f�抿0o��&�ٙk���[=��\� �u`7X����k���_�y'�>N�3�v�x�XH�I�����e����GK�ʿy@/uo�����pj�������'�_)7~ҋ��M*�՞{�-ӱ���������ý�䴁�T��G����(�z�c}����LR�@\�j��TK��LS���/p����������-�:~�w�����I�y�h�A�N,q6]�E�V�]����xt�ˀ��m"�/0]�T���70��5��&]��Y�
�|��&N�.9��Ck�mk�����dT�⦾Zց��Dh�E�ȵ�6�RZB*�+�?:W�vs�q�a<Un<�����0;�/q72��κS�Y��t{��}k!�V�/�k�w�St��$f��6�<> �pE�3�3���h�����Ў����3���Cu�[�����F��7�Gb�{ҀF1O�tmT2RʉM���Y�:�����]����뻯�A-X��?-l�w�[�ͻ"T�$D�+��.^���� ���T�����
����3�`�a\Xf9�=�k���و�^��@�*�Aѿ�	?l4D�_��/A��Al�{��!���ީ������n��Og粙�44B��	�@�3n4���jh�$y�������bi�:vƝZ/f�yw#��{��*?#���PAN�ӟd���KH�2�~5��ݯ��OJB�� C@+m��+�3S_��C�j�)��T���{��9T�=l�s��zK�P��Y�kՋ�����c^`�)��W�����b�]5Yr�C�:1%�6,�Ӗ~*���DC��
D�Y�Hj�o�_��xd���!ڿZW���	�G~s��'��a��I��NP9�'�h{�q:�h09ikg!�Vm@�=_��R���ݛE1�$y�&L�nu�3�=�og3.��A7������}v��kx�	��RL���E�I陏�i�0�X O�� Yr¯��1�¹�%��1�P��.|�}f�)����vZ�~�|�Z����ִ�*v;O�6h�vw�dP��5
���t%:�|ZC_�����80����Z<Y�A��e�zB?x�iwGX�7 B�yS�M�{ib�5�7X�@��}PS�K��U}?��
sd��4-���N������Uv��̼߂\h���A����I爙��N�)���ߓ��+0s>O^�M<��"��9���0�;W���#��фi��9���|�B��"���hL>�2`�E� ��S�A#�ؖ-��J������l�U{�#q
u���ǟ;e�x��A�l֠~9l{=�Um�Q��?a����e�]�͙�S�J��NF��D�O��z.�n(��:X���|�Y�M���>Y>�;f&��Xg�+�K"����O{d�ٱ_C����9�0G�m�H�����0ˮc�'m\K"��H���Z��f�/���j-u��ؠX���F:*o���3�
|J
�*�O5~�H��r
	�=�?Q�[���9$H�Bb�هC&��Tv��Ǳ���T���ֹO��c
�4s����/�fm9��з�F ��k"Ǣh�N��(4N�.�㏯�� ٻ�Dd�)��'�Q^�>^�ItJ}�P�;�^:d����.���m�ԯ��n�+Y�4 �#k�}[a�%Gl�Q�v�q�£�oY�REhc��=�q!r�C�|��[�`��Q�.����q�6Ŏ����o�q�-�O�q�)�3�H(r6���Ab<.�A�_&��z��˅���t���&�jBk�ܴҌ�?/_�v3�1���Wo�tѮh�<Y�zKt[��츽�F�3G�T~�_r��2�F�!)W��Ls�������!eR��c��n���p�:.Fa�S�=�/�K�F� T��#_ـ儼��w3�:)����3�j��L����)	}��"4�m1�:<9ܨ��ѓ)�N����Frz-4�F����J���X���E�}oh92{�N�1(����T\}|�6���K,αj��m����E��FUJ]�hP�A�t�k��{|�\�GP>c]�6���J�F�R��q�@n������c�}�{S�Y��pr���0#@ [Ef�][Ψ���G2ػM-L.�~�S1�u���]^�q���hx���p�nޮ[?�ڰ"�]Z���"\e�Yy;�f��<m�Zv+.uB6<���:6��+cl��Wy�xg�JYde��}�I���x#1���O������#����rb�We��.�=�/�<����U������m ��+�+�\M�@��o'���zųo��Z��19v)�P4��N,{�P~��X�r���c��e��ϫ����c�B^��2�p�I_/����©M��Έw7���ƙ�柜9�w�t�jA�L�o�O�3rm9�M1�-�\��NO&�j��X��oOx�L�o:���e0��U�J��� ��c�����}����{��QVME׮��Z����j~��k�\P7��FUM>�U=���6�H9Bp2kcu�*'����6��ߪ'���|!���av��v`�3��zˉE�P���5���i�Roْ=�	�&��A������#��ڜ_\��a� �j���cg��	%��x&n'ì�'&�O]`b��Sī�]�(
�(6N�c���?c�ާ#�9f�~��k<c�b���2~�b%�����a x���oS�bsŻ�:�!�z7Qǧe�{S]S�u�\a$4�Ӫ䔑fw��=cO�ZU����E����6|���
ob,��Jy�*{1-��}\�ݗ���B0Ҫ|�K��u���/��N�G&�;F���m�/uϫ��� �p���5�;�{8L�,���N�*T5ɢ��C��VE�j
?�������p��t��ޯ��_s3@�a0gR�79s��q0���v��V?��ԏ_@�$U�w����X8��3+����}������$o�V����AN������}Op���j)�g��B��������A]Ǽ�;������)��p�xu��H�~���/�H�:W��N({���(���ۛ��N��Cۻ�N��o}�e1�	D�"}6�(hv�ޯ� \����&�?ͫޜW�ܦxE��N����Y~HF��s�֯���;a�+7��\��Y :C��+rW������I'[�����i#��k�g�E`�QM��
q&:�
4�-a���\%a��i+t"����u�	i��J�h�$l�q�y;ӮwZ�?ڱXе���h�,�U*�� k������0?h�%U��I�|!Q��RT�����3	2��T��ɌšMá-�o\��+z`�'���b�Z��X�0�a�O�ݨ�<mzc��Gne�;c�dF����%��
�,�ыQc緙��5��ˎ����SS�bw�5_���R���7w�)1������,^j|�撡4�i��kۊ�9��1x\�o3O �n�i]Y���	��</��99��ƺ�gbL��(ur&0'�?��#;�9�k7�Qp �A<�x�\��=`R��>���beE]����[�2��)1�>r���.��_�W�ɕJ�| =����ޏG��j�f&d᚞�`���CC�T������8�#��t�V2��T�xv�wt�xX�q�KUE'8`��ܛj����!G�i���&?a���{��i},fm�N����F3(�و�]D�:�Zd�>��{Ã�;�	+rf�_nv7��F�*Z8��Z?S�@GI\��xȃ���`��R�&U��������6�8���O9�����5��%!W'���9 "�����t�	��|*���@W1�ZX�f���en\	W!�����Sl>N��s �t[�����M��T޻;��/a�\O��Z.OȞD<��9��0��U�<9�XR8;h���cI���E2�do	�h���D�� �n3us�ޓN�Q�F��)�I��U�"�����a#�Q5<��
L���I̡�����&a	��2��#���@����p��dt�b��w:Gz���8oº=H�M:ꉸ=�+� Q��!1�5�C��n��\O�0��#��v
��Q��+B���]���4JOy����==O�'U�e �\`b�[Mǻ�O'QK���3���P ^=1�JcxL�ĊQp�?Gd�m�wy��nl<��,1U���Hi���&��eW�m@��<e�l��X�j+38�[zSAB^@(�f�z<�]���L-��\y�{���C����M�����޶�gW�Y�$t��]�J�u��o�C5pvƵ3	����!��YeGu~��
�jά�C�*[�;��@��n��8��*L�fv6�(�st�7��{�R�?\���BܖԜ�f�ޛ�:�.��]Y��5��I�3gRZ~��t��������R�k	�j�8n\��E�نǜkl9�<�8hS����|Y�$%5/p~�X=-�d�M���OjT<  ;�;�Ie���	{�um^� K�x��/2�ᕹ�Xc��ԣ�rbc�q�`�ź�K�*O�M��EI׌�%ݻ����C�bT�	���B�vQEHr�Z�(��J��W�Ai����JE�%r���Y�Q?���!�&�UX#�1 �GWd�ťJ�߫P�����<���v��s�\H�vr�N��Tz$�j�&�7���_l�jdÕz��$& ����ح��q���N�o4U�s�qa�Dx�J<v ������@qo��d��NpN*�}�@��ݨ��s� � �!�D<��f�3L&�0/�U��f+Ф2��*�Վ�P����P�������%)S��ݳ2�N��*��XdJӃ��4Ω��z|�%ȯ.�y�΄[�,�#FJ����v)ԗq��M��*���K���B�?r�b��aE�:��ϼ�4-�Ï��l��6��U�A�.*��4�;tŕ�k\��feKd	��?�R����u���w��L	솨��I�������*��:�� �0M��ÿ/hN�����P��D�B���1՝��x/ɪ~뎃�K�%��8Z�u�X1�&�4�D
�X�Ĺ�S��E�04ST�đi
���� �u!��IS���=)rB���2$p[�758�[�mT��1P�����fQ7�O�C����z0����;�ô��?�H����Z�cĽ �j!�(��8��jTUX3��qj�/mHID��Ӿ�?Y� 8K1��0��d�;� ��a�������;����{�^Y�܆�K����Iԓ;F0�w\mFRj��M����������{�Ԍت!�������
{!/<��,���Ow�}ε�����-�9�5�C�
�>�LK����:��퟼��'U�`y�n�HJu�9�l�nX���zѻ�[qOR��2{ȓhIz�hb�O{�#�{�*{�H��ڍ�l��i���F �S����QHX���l4��D�"b;��3���ح�>-�f��{p��ղ�Qgs#��	ĺّ@�|��[��s���P�h���ȡ8�����P<'Qmv@�+��2O�I�wJ�ЇK� }n�����Ӌb�Dj_ݰ|��x@)�^���j�h]���%$��?�L� �7@�g�����l��;������sM�$&�D������������.�<�N�b�K9�D@d��0��Q�Вs�Q0�Ks����t��t��HمF�
P���Cn=_Hf7������=��@u��)̻	��T�E����:�kR��{���{C�#��H����J�:1��f�������T��b�Ԝ:E� eD0��~�U�4�.v����_����x\0x��HA�x���g���Lħ�b�H���Hl�B�������{x`M�Ԣ]E�Q�X��&T�>X 	�?׵d�+��O�b��5Z`�.=�mW4i�Sh��%y/�_UZ�~4)?�~����")��c���1�`|CD%oS]S��W���n8Í+i����N����-��J�����k4VP��M�H���E��`�z#6l�],�ݔ�ک_�����Ǹ��7����f3 �.+qvY,�ǵ��
�b���Ķ���K���P���b'��j2�@-ľV��-���AF�:l�U#b���+O���z�j=r\5�a�c�|U���kP�ͧ9�O1!B�.RHw��Y�T���r��.($Vp�t`R�wp�l�'"��6�\r��]�/�4e��3�$;NW��8�k��E�hH��嫆,�*��X���bJ�)T���7�������3C�Č;>դ�a�#>-�~����/�������L�@r�LS�Ѥ3Z���-!E|�Wz]�g^��A�ɭ�k�ѓr|1XG��@����rE��L4���n�bQ�;�Da8�H�Dq`d�,?t#D�2�q���Gy˅��P�B"SU#��ъ-��B�
�'b�vK<����A�~'�Y�x���bLM�"�p���4�/0�����*]�^��M��:��WI��Y�����9�|�7n���v����PlZ�	�E�)�����J�خh�!�.����u��@�Ƨ.BU!�&߃�g�=�؀#�����h��뎪��>���*�L����*g#��w�[~G�!�q _�O�{���y��!�#���(��]t��0�Jޱ8����Dy4�� 9�u v�W�$����/�&�w��k���,���"Ƞ��P'~<��	�9X��H�}ha��yɱX��73:�����x=b� �mF�?�y}��F�
@-��#�_IoC������l��`c�����GAZ���[�J�69<�ħ�����	bM/����=�&�pT��(�ina��=L3ڌtU��nr���XЄ8`�[TCSD�x�i��C���zİR� �*��s�l?��EzH`��4v!�=^����|�-�(8��oi�[�>q9�13��ճ�*ԙ��fe�3���!�� ml�&�ˍ��V�Ux+%%�8r@r	�K.�/���v0D;c?Ym�?��b�O��]�-�)��P�T����=��u%��h<���\k���㊍N�̃n�<��M�r��O�:&s;}�g'�_�ܧ��*�2�
�7���'�!�A��m�/fԫ���$e9���X���}1w%�I���1�О���Ze1�ʉw5��?�\D�,��!���.V���W�x��'���m�=���8��ꨶpi$ztQy�2�b�u�j���	�������n H@���Ć�T����?�A&ʙ������YC���Ƌ��W�[�7Χ��Id�i��H��'����
�Jv�_�+�:_т��s�N�W߄���2���箻?ps;�f��˞�_?�iX�{]���
V_�> ���"�]1RBX��|+��h_���Q좦#�eT���#3�����Wa���{�K��
��Ox�����9M�R�@R�.ު$9�L��ؘ���8��1���RO��1�e{b�`T���DM������-�>B):v������.	��T�~��t����.bR����g:h_���M1����J^����oa=;���7e��U�	�A;I���l����������9�x���mΝOgC�h����/�@��i�t�]T'�3�Yp)�E�ʳ���T��=W��0[ݱ��g߸��W�u6��5�Q�xSG�����W~���s����ݎ��ݼ^[�D����e�L���6�مOo�wk\���հ �H�8PE:M%g���^�V�~��n;�ݬL�*C��n�TNb�wL�~]�ޘ��g.�?�E�D��l��XRD?3E���B+�(3���t�w��y�a�
�[����U�x�g�;����sg-d�����B��W[�
~+^���b��}�I�DYH�p����T�,��f���=�+^̈��ln+�rg���s��S���f�u7�&��PnqX%��\�H�_�	�j�[�u*��i��e����*i,���P�O�7��(r�a����AO���)9�&�'N8t�e�}%z.���HUU#����O���8M���7{�q�.d���?~Ζ�r��ju�wy�E�<�t{��Ā�h���9#�I���]��G�;M2J[����S����)�M������+	e6ӹ7�6�i���T����In���	cnߌ�g����z<K���
v{�y�2��5��~t��!�hF,t��vN���xk���}�� ����A4r��n�ޤ�ӗ�~|o?�w*�H�q=���&�hh&��Pf� f>eD_O#����Ԉ��}����ĉ��w�!������ښ��3Sّz�p�a�q�b�j&~5������-����ə��S��h��%��w��0�����0�
��������I	hD?����,玳�N�-�1>�����S�Nhq��ʏ<�-��77|�9"�AvIi[�Ą��6����"|W��z\ko���W�ig��p`�gN�Ee�JͰnL����[%�I��c���݀��2�v�����^RzN/`C�qF}tq���	1bV�]�ճ�2x�2�<��)8Uʢ��ȼ�l�IXe7��D���Y�b��8��;�V����kR���ӑM��|t��� ��ǹ'�<ث�����5zt�K�E��������;_R�-0�;�iD؉ن�Bu1��8��tiLb12D3�bR��q�dh��Z�-��w����ƺ�:���^1D��eK�J��4�j�i��qـ�B.�����A��Н\+�XJ��}tH����&�ﴜ��D�JM�4�Q�#�A�!�Ik_�������Z�ҟX�k��5#(~��V.�=q6��D�X�aR��7�l<.<s���jeg֗j�H]�a��a��S#e�m�����Giq�{��4�gΛ�|��ȧ�8�5�]6�O�H�aN��ե�F�iF����){<�o����'Z\���8<%��L%ݓ�'��G�)J�(ă�NSN���s�kxs����M��2�_�RǦ>O�̊�3G�JC�5^_������7~^��S|�A�����hj|8kب��N_��i�3x�>^�ӕ�<��W�y�2�a��cՀ>�~;u�ߎ�B11��85w�1%�k���z��-.����q��x�@.�7c�}��P�0�����\t�_J,���g������Φ���~���ZCӭ��3�[�$�f$��ˆm��S�2��
	G��g�he�uk�?�.oz�<e��V��Y�f�}�l����Q�r����Z�9�t�ԥC���:5j~/��Li��7��X14���N�U���8K�l�����a�D��^޶�ja�z����Ϩq�Z'�Q������x�0���,^�{��>W1.O�s�3a�;$z.�L{sB[�O�]����Jn_c��D��F��N�c���dn;�s��i �$�]�D��t�3?IMm�5����'�V���:�C�b��u��޳O:��f6��Zd��C��E�*UD����\e���/ic_��#��������W�w�::n�S86����U=�[�`��M����'nz=��;������Ѭɜ�U[Vt�;+�h8*�W���6C/�O�Y�ki��y�)5z��H:7zK@��~����sgL���)YO�<ҽ�
X�7m3҇x�t5b���g�H�r����x��'&AP��ӎ<����TƁ��%�[��v"xؕSy�uiI=%��/�IQ׭���7U��,]�v�_[&�N[�j����F�&�;��]&���}��T�͋�g�r%�^����mf5g���҅�6������p��(�������2z��_Y�45s�7�iތ7)����`)fܙUV�|v��=j�it��v\�C͏oj}_��v��.���Ok�{L�59k3ئ�ڣof&�x�g��y?�Ꜥ�^��qj��.ѣk%����]u�<�ˣ�݌wО�i��%r���܀���	]<�n��GT�~'�'C�}��௉�Y�NcA��p3���l�^�?�G��Tk��Ӗ����i}u�W_��}ȇ{�K/fS[�^Td�����.��gƤq�i)����6���O�ǔ�jA�v����x`��
�F����w��4�׫�L�Au��Z_�TI�[&��{r;����C
B����i�dٴ����CXu��)f!.;vX�n���u�W�a���T
%�A��0B�mmu��A�|R*L�+�흖g7B�QӔ�'v5	&V$�����ĸ���P|Jې��N�9���47ϭ��B�"82i�:z��q�Ln=1��9>pI�ً��A�ͰS1z������#���Ǜ8�P��>x�X�t��t�Ha�Lh� )���#S\ǈ��2�����^Q"�˞��1߷�޼�����	��}�.�Yn���%�^��d��FI9ھZf�ս?�oݟ��1%�(jk����w�sN��Z~�����HuM�!���X;}BB�Ւw�?LBѹ�xV"q���7�.R_&m]�	�z ��J�HC��f��g_�cB�=}�fH,�Y�;nS���`1Z����
��i��Qk�m������`�X|��c)�8RtM��M�D7����qW�6�ԫ��;����d�ѺO��cv�v*�!X�}�����>m���c|���zeǌ����C�Fx`�@��� �3��Rқ�L���O�T 7�e��@�H���j��,%��O���wN�􄑆�[J��ќ��8_�a�vwS[��r�� P�w��O�n$�G�|P90t8:�y�����׽ 8迪�Ć��!���;?��b�
i)���d�Z_����1�r�T�i�pvӴ���/?�@s�[�'󴴟f@Y��4�G���hJC�N� 8��Qn��jd~����0��gM���!�H�6�ޛ�]w�y��7'�#Q�J㾗~�U+cf�|5`�Dt��nN���0�� ��j������@h	܉>�2��{�ĝO���c�-���k�Pa���� 5w��B���9����ѓxG"����a�~�l����X5�Zp���>�$���'�b�w� �~�5��w�^�72N���r��,�L{g�� �Z��z�%�N;Ih+��M,��5��ZE27�B��͕I�hH/"��9���t}��b��РbJ�y�'�A�ɣ\эJ"em$�'��!+Ox�D�+�x#���m�zQ⸷���i�Lþ���<��~�0��U����P�*q�+M�o���*gAOM<mکA�Fm
�m
GZQ����}���#��=1u/B�x:�L���?��)I��CYA�Z��:�쾮����9.�Ȅ��x��U�iڊ�R	�|�$��:� ���O�6]xo�߸�Ï�|F�SYF}��w&�Į�7�N����XW?�&����-���w�}|�9!:5tLc�˭�4�3:�DY�X�OSs���d�z8�(����@�~Y��HiL2D�j΢%��b��΋�I[$<Ɠ����r f�o���M$����bD���Py�����C�r�x
���ף�� O�~/mJ���E�'����@;����-��jmN�į�B(aH���V�2ӵ�Z �:�a48���c+n���!�d�n���WD�_�E>�-K���S�-�:Ϛ��-�����	��(1��y�S����bP[sZ�}"�Cщ"��wL ��w(�`�0��o�~q�L1~e�z�����i�𴓎"��(n^��%�S'��_�<A����\�Ͻy��?Ag�ヱD�A9�^S�G�:Ju����RPұ=غ/�/L�s�����L��4�CM��� E��ɧ��������K�o���PDhHޠ�'��|��Rb�}�{,8�~s�wG~��g��Vd� �nRp".j�麙�ŷm�L��ks���������o�)_�t�f4Ppx��O�D�=]�f���K�H�1;�b
�y�|@b*����r�Y�w��\��������!)�Qu�PU��Cż��:�K���:k�?a᠂�
Q������m��[�^������oy%^��ﾚ�Šzg�h�_'�����b�-� �y9��,��o�[�͖H����l�·#-A�ߦ7i��9H� KE�hj|��?/�?H�]���x ����{��i�Sa̋��_!����J�R�߄��3�(�/�%�
dI�f��/1h�3���
'�^�b��1���L=��S�C�Z��L�-@]�F�o��݀S��8EmJ��r�nҳ����lZ��B���1y�cXM���A��qn�D6
O�CK���䥶A�]t�;������߇*m�"�lz���ܥ�/)��׋�r
DU�� _|{��?j�7P��+7Cf􀄅�HT�]����4��~�qM�|R���2
�����P�� �-�zu�3�a��х;�y���-z�M����QP}��Eڀ'�������$;G�d�_�X��A�߰V�f���U�Η������2�.P:
*�;�%��I�˨٥i��bZ��X�Vޠz_�r�K��6��1ZY,}�#�H����c��]w�3����	R���/5s���?�Ca���6�b���%^9~^.Jغ���-��K��1*C��r�'��?��d�|O�����G�K)�F�'t�S��ρ#-�ߜ�!{���9��ȇ��(n�)WE9�6d Q��"!�w���ŏ��!�Rɞ�~u��qv�¿�Wr~�^�?n��X�4����Mƙ0�D��Ma��죋���p&5w�Z>^X����.�

P�����Re�j,�;ӘX��`�1\M�l�p�ͥ1ʙ�q��czm��T,]���$z�F�tN�>�η����R�]_���/�1��fw�\xUzTN󕓩4�=��Si�2�>�L�E��  �$j�Z\\d�kpL�S)��5�G��&q��%*Ei*H�<xme��+���vI]����Ћ
��n�D!,���|���X�XX3�vo@s-�׉����s�7������C�D@�H�
[?�G�giP�Y�yq���Przs�������M��:N��2�`�b%p�_�`�1����P����^�.�uH?�����_͍n����Qvs�m����HeJm�<Ԓ���W��y&��*���XH5��x*s�:�v ��u/�� ���BA�f�ț��H>&���"�\�[��6C�4�_:�8�mn���"C�8�V�C鞎�AG����E�dSp�sl$j"�X7p����X�!�u�W4j0���SƋ�C�t�j/pHã/���'P���?~gR/���#(�τKǻY&{���9�C�(7��_W��-NB]f.�X���O�4�ƧF�,�	�#C�	�>���Ρ%5�6ɋ���.�_r��K�6W�6�8*�ӏ�[��c�&��UK�'��y�]H,�� zb��;��b�a}[�ԜG-p�z]��~fڜa7e;�C{q&���s=7�-7�]��ҷ�g\�
ϗ��hR |�0����#��6�A:�Љ��#f��YɊGޝi���>.YB*h�g&�vX���D�
7�3��+�q��)����y'$)�4�{�E����`L�Ʒ���26;����R[��� ��Y��C�ݣ����RB@��v-p��:{*�4���_����ct�K�-q;��Kw�UA�D���ʎ4}�?�� [9)(j�JI�	 !`�.��i4���MJ~
�/-�����e����;`�f}�@|�Jm/{� �]��Y�H?��7��q�  H���־���7�H�R�Q#��.�ɲ���2G�=�z�ͦԽ:�/�@?��\B�~�j[W�Tж�$�3dnKpϦ�RNH2��¥~�TS�q6�>9}g��;9c��浲{u��3�c��l��)�P�s�~>7�J�͜�-O�z����{���\.�&�kw2y�����/��*8�?��>���G��?l���t��G���6�D���N��~H�����<���oKCy�5�9ͶMu9j#&H��6�FU���Q;\���(^�>+�-������i?�B+Ruͧ�I���X�n/�e���\�k9U.�yin{]3��d����D<opl5<-<��/$K���'y
��-��_@|��vU+��-�<,t�v����{��454TO��+��։#�Ɯ ��'���5�C;����(�*�v
	U��_p�/^F�Թqk$��
e����q����/3 eD�9���f���d:vZ��m���;R���}�]^�9դ�^Ȥ�5Ri�r?{�#�jؘgj��X�ˁpT3{5��|z�H��qenZS/�9���$ˁz6M�pL��ܸ���nB�\����N5,q����V�][q�vu%8;{���%d����bi�����^�J����ڋ��~(4Խ�x)�2�J�quLm��v�)Ԉ��`��^>��
�w�;��m�d�t-8S&�~�n�Ƀ5��E�>"? �?���%je�Ԗ��:'�$dHW��Q�N��>�:�O���C_�xb8Y�n,�q/m_Jb4��>1����R��W�n�ժ�N�4���[�p��<_.|���_I1N�zҨ�����-�UW#���Dee;����\�s��`m�B�������yt��qm����6�
YөaW�N8⹌�nj<|�ʧ�M��T�.z���Aw�n٩S��Q����V�G�V0�n��»�����d���T�i{"�;��ߺ�t��b�͌#�i�Ƴ�ۺ̞�H�� Vn洞��R�K&����ǃ���MU
+ٛ�D܃�o� �K"�)�c��4e�<%��p�UUd�Z8b�:�1�%���<c�[#��������G���<c���ItB���E�*�u�����+'\ E��磞�V1���.q0����=x�ў�����og5�yױe����[�:�iI�9�$��)���(�ˍ��~�v�9dB*j��v\S��C�⪇+ﺪj��ƕmn,�$#G�y�� � 4.�m����0�sa�2RvPU�X�k����<�����:G?�p�����<=��<�k�<�87�������ҫ1�@Ч+���v{��ԧJ&�{�y-���[�[�׻^;��%�X��~�s���U������\k(^���O�+)Ó�����J	6�0�EՃ�I]/��o��z�	�4�v��u��~�#Ovq��?�y���j|�S%M�;Ŷ��9uD����1]BjjaV�sB��(y�!G����x�0{��j#�� {�m�O��nt*���B�˼S�5������p���L�WӦ	��"�r6��"4x�����������J=���)��T���Z(2aZP�ٙ�J�Ǟ�bHJY�T�^dO�=��;�w������>��|�����?�Ϲ3w�E����s~��$H?t���b����3p͠[�C|�R�n&����ϗrf����#����֤�Y�'k>�t[	E�i�;k����{o���z̶���LG�zx��3�`3mQP�g���(kFڟPQ��{�=l����E����uLav�����w��=E|�\���0>�V��]��� t�>�i|RQilŸu^��M��� 3��5���H����W�Z$]���#�{:����a�_��.�S�[��'�L��� � �ׅ���t��^7/�P6f��Q����|�Z�	�/-/zn�N�y6�a!���`�%���}N�
��]x0�ňP	���M˛���~����ԭ�bD��|�����/"�#>�[S��7�I7��v��l����l�^�d�?`���J��E��S�Лα#f��y{ 8(��	�_�,�]�B�F�۶B��c��+�ߌ�?����<h���z��
�u��}~�&�nI^���L�٣U���ߚ�����s��RS�I]���{'ނ�K���җ�i�+�A����z��Y�:��C�����	%��w�K��kv����h�0��	T0�K�\ҳ	 ]R���)���ۈ��P82���#\o��Ex�m��2��z��9SajT��_I��m�B��js{��б�[�?�����C@y>?hzlb��g�U8y=]�T�~��<��	���u��B$���\�J��,�gb-�y��0'o�j���O�$�Љ��~�u� X������'՘���|����'�г�b+�XhD�)�ʯ|QZ`�Y�� K딓�6S`���LJ�z4��Lw�8�i�XRC�yQ�Ά�l����K?���c+;#�$��y��A �b��P��0%%����������AI����ATsQR�&A���K�[���
 ��S�EW����l�ተ���:�Az����aM�b�����^Iv�У�t"��&}��X1��o\�Dd׽A~P������QK�xE��G q9�6!�+��V<~����&%�#��S��<�0���a��6�]i �`2��2P.��Y��j{�I%F���Byվ���]���͔8 H��lR@ki�y�y�!󋜚C-��V��t���>�e|VR�yh˹R�x���w#"���<��<�����v��7�$hӍTr>y�_R�t�?hn�iܫ
,�F��5�q�4�V�l�Ƣ.�U&+��Y-AZ�7��F:���6�_��c^1��u*J�x�z���V�<M��
�������!�S����Ψ���/!`\u.,9��`�h_����_�";�K�}D�|��E~XNe�ê&�������T�������a�N�-�P��v_R\N��ܟ���e���
R�r�DHG`&�oJ6u;tTt�=�&��+�Η�@��}μ �g|wV�3��5��x�����*P��¼���2�%)3VC_������+ѹ�AMKa���s���2t��7Yee-��f�և_�bL'~�SB���ڒW~�*�[�`i9�qL����ҍu�b@�;g�j���#��쮈1;(���-lc�8)������\�N�aj0�OJjKYH�\�B_UXL�Á��ϧw��r���N���r�=�(("�u��k(Dm��b�K��N�@m'*m]EY��TUk�\�?^ԕb�?��X�{�R���+�FX�K�Sk 3q]�?D���`��T.l'@Y�dc�q����<4���m]�=]�+�Ʋ��FV	+��\lx��3������l��$~��4�I��@�l����b^N~Ԇ��1,�z�W���1Y�hl�j�Y����E�:�V���y��?��	���-F�y�A�4�<޺3�ﳟ��W	�^5^��;��`�l`�Y�	���?������y��ZE�9c�)-<�f~�c\8]���$|SE$�\�>k��#���PU3����Q�n����������A�S��BcQVh��I~�3^�4��5b|Z�~ �\c! <�e���p���R�������C�O�~�9IM�0_*+��u\���������"�YյH�!u5Ξ6E�|�Fb����"Ҙ��{���%Q7��ձa��VBmL�ɔ��MCT�0U���:�2|m��' ��%1c� ˵+>/���ޛ�eU�1���vv�T8��A^��P:#`���N ^�R�*�$� ��?ő�]���/ރ«��g:�[�u���sm>8 6 �Vt�"��>|
\��&����l���m���� ���U�ٷ��Yl��2��P��J�٥�nE�*��ف���	xRb&�.�@З�/�
qs�cR��H�f��������V��F[f�.m��'�C�1�m}syq����d�*X�y}�n�=v(����ї�	*�+Ũo�,�G���
�U��Q|D>�_�{Q�x�1V�#�Gٰ[R[��]!�����<�o�y���&�y��K��o!tN�=3�W�,�]��G�������|�*�����,]�equ�����WvhK2�8��U������ma���9Kګ��g�m��̍����DWn�J��f���0)��\�S�mR�u�b٢���v��L.�,}�X�`��_T\;�:�`�X���%M@T�Z<^U���5�&~�\���@�F�*{��nK%Fv��7���1EڻO�KP��7QA������4�ڬ��u��>׌�L�BM;c�5��|Y��Ľ���S�F|!�"g���@ꥩP5��3�vn������ro�g��,L�,9�DD��l���>�}�i"��Ce��N���٪�}��VPJ3�A<ѭY���ߩ]�	�����F��l�oG��w�i4���x�*��`�!I�V2��Ï��i&�5�|�g1�t�5]��3v\=�#�c�����@��ύ�E��hV��sޭ̸�g�nWqWūY"3)m�qm}���*�0k[��lB���1��=]i�*)���|)�Fti���Y�����{s����H:�ژ���l���/�3�L�����ըx"�
�?c��V������_��psd�uy$%�׫�W!���)Lm��C�s$%ň��}�q��<z��y�^��(L1zl�r�ӕ�� ���ۏ=%U@�9����m�הּo:��$�Ի�����W��uд�����a�`Dy���,|��8����M��*��cIW�0��.D
��r��"��Ct]n�<ba��cq���8�1m�yܭ7�L<�C��2�d���(�@�ׅ]�In��f7r���V�+v<\�$H'��0�י�[|�_�/�z��78�#���=^�T��ű�aˈ�r���Oa
-\�1��S�=�7Mu�N]$t��M��n�K�]E���̂����C V�o-t-wFg��\ي���I&�c�m���=fl��A�|;���/��ʰx�̈́�+�G(zDZ����Ʈ�!��Kym���G�7��%�"J��lw�����^�,Z(�ME�	���c/]J��I�DX��:p6�p"^}�[��U����a?�����u�[*��.�+��L�/6��ի@q_C���N�`����=J�7�_r�j��j��̎�c�:�������Jj���N���"n���;�����v.F�K���FW|<��K�W���H�}��:���� V�����&����HXGRd��-���m�0_���HXF�)�f�M����kI1�J]��;�w���u��T,ў��n Ԓa*��! ��7��:Y�ԧ>s�-�u Z�+��n�*>nn����v��	 d�%��K�h��ߦ.�l�t��#g�I%���*C�э�f˖��4�y�6��iE�ϡ��w�^	cB��C�V��O�ˋEm�9��� �7��t�>����9�u�����A�Ins}g��������`�С�R�8�&p�҈p��qхhw[?t��io$-�I ��W�JxlB:~�>��oj��~��6� 2T����O}��++�6�����m籟21��U?�Բj a�^ځP�\"�Ah���&�_��*��u�\��f���=�79��b�W�T��֠�S\���_��]h_������b !��8��j�@�Yӷwƺ.qx���;@h�G�Z(X�NcTI�l{\2�@�4t1?��y}��y��@�Dn������N�I[�7�i���h�z���/GPO�cߜÉj��HSI1���,�^�
�ng�E[Q/�ڴ��ϻ]�[����'�Ae!�{������nQ����w��iIc��F6�gj�H%��Hsݐ��ב���> �2 ���!�:�FR�Z��2?����C�Ŗ��� �>�K�G"�G�$�;�����hg��lz�]�d�b�]�6a����c��KK㖋�Αˇ�E�j�[�c�!��߄����Z��ŲZ���FƳ���H�OױE�#F����b����}�_9G;Ń󇾚�Q��ߚ@�IY��mU �2����yhK+�!0�mv*c���e�����A�?���!����Nי-�_2���cCҀ�{w�����+�ed��FI_�B2}ض8�{Bj�)��.OVIB�=W�gO�5�A�L���o�vL��/D��n�c��t2��^Vk�E=I�n��nש(6um�h�/z���>B	2"�@�,Tpr�\c�#��ʰW���$zt*��Qנ�lfatO��7��&���G��gl��|���M����pb�h�Q N2-M^B[��T<��KP���B_?����y,�t@��s����+��	��P�<���j^0��#Bv���_!���ā˂��K�Ϡ{�a�M�Y!g��=�L�ʼ�3_����& �m�}#�6��,&@2��*˘?�����-��2b�Q�HghI � @^V�j���D@���ר�)���_�Z]mD p������ ��sϰ4��µ�����+�s��h�/pr�)zч��1RXɎ�p��KV��^+�"�;���ا0�ǆ�n�p� H��c]r1���i~�T6{�Ģ����☖u�j+#��[H�aç�OH��譢x�\d���Ø�|^����<M����u���s��r�}��~�[ƾ`�E�Cf������k3v�*�z�t�5������J|�#w��b��W�4���>�g�3���w6b���}P�Of�������mOqX]a�^�o	4�`�⤹/J#&���@F��:	Ҧ��Hv]{ꂲ�M�����0�s0�?�ȓ�nX�ex�>�E�j��Ȳ���ai��=���t��/�Q�A.~PY ��i��3�FK����j�a?��r6G�FE�lފ1�����'��n��>�Z�e�LVB��������Fg1\weɶ��RY�6�L=�6��ʖ�D<F��Ff=�  T��Ā�#�@����/z�z���T͏���^�V!g	��̋��d��~�"1�np�x�q2hH���ԩ�_��i�$F*��όD|NWx�<�Ѯ�(�L⃘��F��񣚄��64����r懗�W�
�:	����- ��<2�i��14��[��� ��~^�Mo ���@��O���1�_�|SaO���Q�����n�*HRؤHS��ѕ� �G�[(��]u�E?�컼���:�?z8����.H���הF�ɕ?ڷ%Z�]���d�`�N\&�`�&��ғD�Z�FP��ʵz�����W�t��!/یZJh˯��+cL	�+{-�]9Ni�������!�v�./��
D��T�����a��@h&�ۦ�`j`I��z���%�7f�&z�k�b)���}��| L�H��ň��-�Jl��x�LIf̧��'z*Ǐ�.z�����?1�C�o��>�5�3�4�E|Dq��{�Y�C*��d^����*�F��d�		�%#���\��J�Eñ	G�?R�g=]����%�����ư�L&���!1����spf̷��|�^�m���C���c�^2[F�VF"%{�9#��)'��9#��h���/���PE�vn@��t����_4+�W�sd�)���M���G�	-4�Z��í�;{��l8�щ΀������~ʄcZ�݃\f��c�ܠ�]� �lBtY�^�1���C{�{�2�3�.��j���jYۊ�+=��!�/A;GS*��*��Cdf��he27��yx���2�Z�6���k�G�g�Г��x��Ht:}+u��ؤ�/3��49+�Q��V�ѥ	�� tR1�0?{BF�|~��̮�w/-}_F:�6�����Fڏ�R�=�pD�7�����n��=&X�r��G���B.F�`Y}r��K�v0oy��fgg�FR�;?O��Z,���Z4����e��6��q'��-M�7,�H�?�+�
H����{1Y}�z�o(5�׉��~�XB�Z�j���y��x��2Ԁ��P>Kq]��_ rG���t��xp�_v���d�5t4p���M�[�(+�����]�F?m���6y-����	�R.}�˷����(��6��zKz�� 鮂�<Pu5+�=)�ȱ���X�O�/Ͻ��8؝��67�+�s�`h����ݎ����#�Y�@��3���zt�\Ͽ�3v��_��~��[��%���@U��<%�ީՖ�衡�X���H����	$-+&��1<Z�I1 $��s�m�M"y�L}�����R	7	�_��2���+�yy����	�
8C��h0��b�?� 擲�b(̗Z��
P�YEq�!ꀂ���������G���&������,���XVAb���t�c k���H�5}��c�!�>o��@��Bep���E:��@ɿ����S��>���Q�4 �H�z2蟕�;��V�!�ד߭����B��Ձ�r��ͪ��W�@�|N�y��Xt�#P�y�J��Ϊ����D��\�#4�|t����F_T?Ot��̅�k �ߕ�)���dI���'�V� X_T|���2.@��iڎEר�����a����EK�3 �!ତ4�+�uk�Ľe8���{��֙���#��V0d� d�]�����t${Z��:���^MEU�[�8un���Xs:�Ջ��*.�Ry�"c���}3�����?`Tb�K⟦�!�҅��x's�c�RoH��.jI��,��V����iԭVA�u��n(�=.2k�2�\�:T%<� ����|������q���]�Kn
5���|uR��������!�X�Jg߳��"[�󬚽|���]Z��p#�z�.���ֻ'fe������7~�#I?�*/�0l�$I�s�G*sZ�ж|�/�mz����w�Tۍ��3�@P�*�q���|���f�h�1�_��RCR���d�ze�~��f�̣��y]I9<a�zX�][�gq28�m���FP1��5��>�W\��O����o�߮'ޏ0_Z���e�m�I8=TV�9���|��X��O��=��s�삋'������6vL����w����f�]�Y�P���e�vS�'ob���+4��u7N���uZHɡ]�� ��0XX�Ǡ���,�ʙn5}K�;,��M'|�.ZD7���l>�K��+���45���Ռ�.EU-D��!���ϟ�Ħ������h��u�<km'~��W�g�_b�r(v�uZt��歺��D��!W!Ϲ��*��ے9�W��f���G�q�!��z,�~��~�k�_�o�v�2���*x�^�Un1��\A
<p�Au�O��&�1!��]��!)�̙�s8$1�Z���˗���E!��_A��ӧx:�?,q7R����g�Cٗ�!��5�����{aR�e֢!v ��>'�:窫p\}�6�Y�$�hP���L�/�Q���r�쁬(��i���(�e݀/{[ߧ���6��2-�9�.�@�8��l6t?��TM�.?��|�yb���بݜ�'��:�e+�i���o�O^���(�h�'dP����6?�Yup����l�%�v���<��ݚF�K�}C#����0L��)؊1�ְ��2�t�!��3���n[�Rt��P����x�U���(�-�����F�Žߩ��@�.�DbT�=���R[�(b ����G�g+�� rd�A�6bʿ��#��sd[Y��p����@��^(s�ݰ���';����ӕ7i���Z&]��e����c6�L�!L�7�c.yu|�K�_
�IpO8;H�&w�RR��]u���.i@l|{��^�l�Wb�ǝ �*Jxա�=S�> ��:-�Hd|�A�пX���,���S�n�u��A���uT�"u�(&z(q�?~nz�,��|�`�⠽eXU ����w�,�x�G7������c�`Q8����|���huQ���g��i�8��o��� Ф`�ԋc6[�����&�l>C�����&�\�ͼ<rIg��qK���u���c�=U�]W�θ�������X0.���Wn�t��ݜ��(���z�����c�K��:� �������}��^�q��W�q�$�+ƽ�֨�OkM��i5��F ���g8�޼}�0��9=пZ�Cj���;i��������)-����� �$~�H�)�-tBr+ Y��̟��3��1v�0��i#�Q8���[�7��F���o�V�cA#}�����e�6�.�4E�X�� ?��1�MwD����d�O�]�^[(�����[�+����Zb$�S���q*�˽=j�(A{P۹F�v��Xi�,�c��ҡ c�f�^��ÍP�W8�im$5���2��rԄ��rY�(���A�胚Ex0�=fC�����2��¢�*�@*SD��ǴjE�Z�`��W6pV�N֫�-��~@��,y����i�U��W�4�fg|���E��a7#A�6���3��ǚ�c�u�q(��sh�F ��x����j0���5�9��|�ҵF��o��@z5x7'�� ��߀K7���[8E���S��r�%�cV����UK��s�����/��޼��r{���`��i�s�(�n
OԖןb��-e,��^
Dmp�1��؄r�j��=Ke���r6̨�wXy�%����8�9cQ+M�� a��@�����!����� MB��0�3�n@�� �������\L4���O���	� `�L#j�oO�s������1�X�clP�
�~���j�� v�x�R����oe�{���YQ�{1��-� Ye��N�O�)�F`�O,?�~�����sg�².D� 3���Qmr4p5�!5��dX�Ӥָ�F��N��%b��;��jB�h�;Z_ؽ;J5@���];ʃ�iR�5��@W�X��Z��^��j��W�c�é"j�G��9 ��2Şog�.�J����l���0)�P�r- Q���X���XH櫿?���&��P�V�RV�4fz�>KY[Y�Pbݺ�"�Ŷ��"�|e�8��o��
x2��
~H�4�!3k��ӣ�Ig��c���.̽�-Z
Ar`k����OB��-Ɨ�����c��f�3~�̻���(�墱�k:Q������&
+.:�?���-C�CGD�7�1Q�7]�Ӿ`���m�h�$a���Z*�xr.�d��
�|r�O��̸�tb�������:w�[p~ ��|�	������B�n��R���F��?�,M�حE/���|�h�7��A�e��٭�_�Q�#6�{�+���D�}��l:&�_8M����� ��y�}enڃFY �liU�~q��򩧫O߈;��r������Kο�pC��kL_V���Ő�8�p�3�3a�gZ�g����4����y�:Y�U%�E�7]{�ia�5E�c��y�_Z��D��w�ȳ�@�|�^���Z�M���S^�h�ݥ�|%�����c{E�S�_�[^RC ��(�,h@j8�����5��X�g�' P���qʓ�˞���Q� ��Tw��\�N�%K���~�E�6��c� �.��{������j*�G&ت ج�����d���1S9ț+��9e*�9<�.�,�N�ݥ���+;o��(��e�|r�y�L&v=g�f顆��]�-K(ڂ�*S��SB����}?�1�
`�z���bI��R�!ȑ��8q�HX285�SC;KV8�%`�9���qdl����5���J��+`�M=ʳ��/������=�Fˏ�����%�<	�*2���x���[��b����O*:	�C����m�%�4![�;����-�0Xt��P�iE�4[
H����L�}�{,��~�!n�5(�җ���aO���Г����$�
�!;��U�\��e�N`���Z���'� ���:�,�!�zNw�_��<��>&X�:> �;�4�N��}>��~��Is_���/|t�1��{�<��W��p�*������vtk,t�x���]�c�f�;��y��1O��@�'��-�8���-c����*�oG��4���M
���>FЇ�� �K�h ��a��%���7r,BZ�K}~0 ��z�$0?��q�_ve�94Z��X����+�^�	���3rB��z��;n�V˼���'f�&�&�m�����3K�7�i6�ԝ����������h��,�LY�w��dA���N:Qg?�`2O$�H����M���A��N����0��:���g�P��V-��6��i�u�0�����T.�AǗbHf�{�a&��Џ5��kӋ_z�%: Ё�������}Q違1��˳���d�p&n���(�<3����B����gԯ��՘�Eۣ��O&z�M�4����f�p&c�dcy]�T0Vy��!@i�MF_�Ͱ!�2	*Y���+΃V>�F0����'�5��:Fa����5�7z|v��B0ܩ��7���6�X�=զ���F� `h��o�T�[�(�~m~�L�߳=��;`<�\%E���-@� U�(�O@C��~��S�?�`�B��??6R3��6 �;���$Ւ�߶u>*���W�k���S��ZD�c��:��"*�SUI5��)m���3O ��;��AR��װsz���1 �T���K�C=��9Mb�ƅ���|=�c�;��y�{5�<�~v�/�� ��O������@���n����3� 3�
D�o�}	�0p]@]o}c�1$��Έ	�򠁜gҕ�
���X�j�s�5�H��e�s�Y����`���r1:���m���:��������'p0Oa�ߕw+ ��_���C�#_amZ�6������쵹I��~��اiȶ�
 �\�*o��g�[w�Z�9�,���_XII�B��l�T$���JnLZ��rꡣ8R�d��:�[� ��a���Pf� ձ��_4�$�<`֬:�aC[,cqp?g��p�Ij��}�SC0��Q_����z�� �������>���N�n�/���?���%��W��/��|!VT!VH���½p�s�F W6�����x�/ڋ�����
_��Tg~��,�w�Mx$���3��<��Q�k������8i?$Kʱt^�`�;cM���1� ��P�bS����W�)`�l����1T� W�f]T�1���@�m��x�g�5����U�(T�g z(�/z����X�Z��B=e=ق�D�z����S/�2n�j3��YM �yβn�ڹ�C��t�(z��	ڝ_�mcX~��Ƽ��-�@ka������&���ԇbG�������6��X%i}G�q��D6+I�s��H|�z��H�ʃ
?�_
��	�1� �^�v'wn6Ⱥ�ȯ�����
�� ڳb�AI�Nz�/������?Agx���40�UI�d�z���Q�XzȨL��X�:����=�Ҩ� pe�t���� �{���`����<��4��:�[7�)�����9�XhcWYQ8L�l ~�K�������$u����6���A�o>�K�� j��7(X�*�7�cUy�pz$ik�~��h�U_��T����~B����{D2 ��+ޛj��= �lNwmv�J���9��Qu�Q��e�	�eDjw����w�-�;6�+�Yk�u�0"<�I�D>`����rF~M���C)u��,���]u���<��[
����R2�L�U_��j�i�~gbp�e|��Y�]�֝`6|K6��/��A�TT��y��,n��
���|� P�.)α����/��Oy��l��`#�`#cP��׏�5t#�`τ^��p�_4m���[^f�Μ�i�i{�wC�>����&&�u�gI��?�J#���nݸmn�%T�@��s������H����Ot{w���<�OO �������&H!�=�˸}e��g.f�æ{4�����>��(�B�D}�����[��9�P7d�X y���/���
+��~냖� ��I����A�e����]̝����0���s�[�3u��У�B_n�]_d����R�l��,D��A�1zQ�9�\\7��cqN�<�O�ap�o�����_�ǻ���g*.�,Ԉ;Ŋ�| �𾈑�^�P��)]��g������Z��6su2.����i���DocK
�(��}��.�� �����@���^+e�o{G^��WaVfC�e^��i
-L!Hhv2lp��r�@>+��(2�I����!����-�!ӡ�I˩��L�Za������h��\�}�sW),֪A��Ș��-<�bR���U�)v�G�hw=s�]��Wt�T������A�~��Tť5���%�Hk��-�<���D��p�
2#�C�l@�5�J}v�z\�@�íY���kP>�����W�����}�v��3z������	0�"�<�"���i&R���ޔ��[&5RAeZ����;�9u	7��9�GF�[�P>+>A�-��sR�5"�_���PuO®Wo[�+]��;e��J�%!ƭ����ҵ�4�����"_���H	�������*�OL����^��&��x�<o�1u�/��}6��9����Ow��52�?���[��jc\<g�c��T )VG�J�B��~i+�ֻ3��{z��3�,��� �(u�Y�-�����F�wN�K�l�Q�m���H��ڂ���
���`���B�+O�Z�y��M��5�(c�D&���5S�t��CX�ӵz�þ�L���\���Y�26�S+M���uܰn�m�'��Xt{�����7��V6���:�Ţ���neo�����,��/j���ک}���>c[�ݴ�}�mE7v��'V��E��߹��*]8s�yI���]8����LsFS`zN� ��mWĐ��4|u�u�J�;�����-r�I�����CF<Y�qqN:���`��Q&~�)��-�k��h؄���I���yv��aL��T#�wh��ja������fY��C�>�)�XL�u���{A���:SA��ݖ��敜�=�;o{¯d�ߒs�]�kF~>������Mm��L'�3����,�:^�ZvU�5���-����PE
F9�-��|H���i�]���.��A�$�*�ete_EEt[<D�Yi
#]��}�	���T��}|LS�V3�ON�O�e9)˂���3��=hv';G�}J�imΝ\�<8J��]�~7��Ott��ʉ`W���I���g��Ԛ3v���ݳ��=F����AyH�ͺJ���_�tPqw���[��x%FȌ��aWG����:��?|{���ǉKrI0�����?��Xfv��
ל�K����v��<&�9�c2�0��M�17��	q�5o��$ i����x(���V�X��TS�1�퀟-��y�鋖��^��PI4C_�]���S�����Y���I�ia�gn�5%R��{�Xf~>�	�g74�~LMy��ven����V��� S%_4���)O�j�r
�Wv3�H��c-�����Z~D�{x������N"�6��OM�`��l��I�e��">���I|�՜�}_�y����s�f�nc-iTQ�w�T��U@�2l7m~��U�SA��5l��=��7x̬���Ύ�	c��G_Alș����A,{������Э:���|�Q�K׹C�]	���X ������ph�J�= ����Y�'�7��`�A���L�>Sģaj�����d*()y��Y�X�ucn��|�־��9���K|���N��.���{��4!lm�')��K�r��4�.�j�oi�!/����}G��Z��IG�q�_�x�M�*�/�#@��R��M��ח8��_(_f鎛���#Տ��4ݰӁ�@�*<-�+9z&�N�D0�0[=���ЁCY��s�oMenb݀䜓.����Ǻ%Q�ĥM��$���H�:J@(a-��D�ʺ�� ����ݢp�z��dVs�bhO�{���x��r;����z��}n��Y��ݕ���霫��b:��k����&���8og�������~���z6d�?,!��t�� 5�*���*��X�=$�a��c��O?����)��W� Nz��|���[*�kf��ao]wAڟ����hW�w��4G��ץ����������Mi��x�4t��Ȫ��a�Ks)�����ebG'�:U�_�ퟗ�*_���n?��u1��Y����[s��=��d��e��GG
�뺃2ޒ>�l�M/WE�����q ��uͷbt�<񝉉2�^w�V٩��I�E����'��S��� �M�x���_v=<�EK�����_�O��P���_#�|�=}k���]C�7���ux�S��g����S�M�x8x>ms�%4��F���k*��Y4�}��H�AP�v��O��v��~F0�(��3�{e��7��m��f��wW��'ؑ�`�!Jn�gzI���2� �Ybcz��W�|A�х�4��=�����
cH�.�?X�n���!��ۻ���Y�tٺxж38W�C�R�uKhI����x��uKe����o+�z&�3��� �+HďI]��D^�PR��[�� oP���٦^�0I���<-�]��������-8�3�`��� g2��Ot���/�#�(����x�Ľ_F\�wFʳ\����Nl�1N�s%������V�"�r�n=V�{���{�Xw0��X��T�b*������|��EN�_�A�D�?녰|]Qz*>����'?���]�:G@����7y��6C�����a=4Cv��Tj�?k��y41�?;܋���m��<�ޱ��}zc�Q+g���{�Y������|�����B����W���a��@�Y#�_¢����0�r�dAh��i�����C��Hr$�~��DHJ��S����	qA�	�Y�8Wc��Q�,|��y٠Ox�7	�����:vnB��s73J��7��pZ2JM
ċ����3��*��NH�2?ϵwZ�³묓��!XE�7c��1���\{X��,�'QC���8&ޮk�;�z4 x.3fw�&vK��4����86�0�Yҥ�)�0�	������_��ڋa��ǟx�1&��G��	�\��0k���#nq������׵�ʵ�գS4��˗���g�'[7k��8�XF�B�7��G������i/�P�ƪ7zE�j�X�7�_ �d�[=�����&��J�^P�(k6'������ņv+A�OH�Z��C����i��<"g��R��v�SO�WRQ���&6�.t֞��I<5�O�X3<��h�-���Pǉ��4���;K�Ӻ��U�����cSk~e9�����H���AI�B�E��]$�VU��[���������Uż����y1�)=�m�����ݳm�j<��<5�2M�?<�� ���7�ߢFrϓ[����(�'�җ�q�ߦ �A�뺆jQ(pΈު*{8q;��H�^��$�:�q>���8v�sJL���
ZxW��?�[��H��@��f?���NB�T��+ƛdP�
 �d@�����{G��P�)؞�f�z�u��?_k��t��o��6x��P �v��,��ފԇC=�����)��RB�r��P��G�.��Kś吞��{è
��ph�v�f�O�\����@�*�g��c���`�4 ���]+�3pi\�#TW�[�w&_�� �5��H��؇x�=�H��;DiM%Ep��l�b��4�3u���w؍�j�سН~�]/:��:�t�ǒ&u�>Φ�NR��T���c{�\�?��	f>�D������jΚ����CB*��D��M����|Q|���.�'��'��ӤQ�m�)q�����G��l��'�UJΗ՜4�tu�h(^b{�����|�J�@��B�j����ZW�oZ �<J��O�z�<#����;����;
b�CI4�F@��t/O`��ˣ<]�Pah��r%�t�qA��Drz_0LP7.����u�ۺ����ӣl�@{ʚHmw�6m�����yS\��:��:3��v��b���}i�dѯ8��)7T�3�v�!y:j��"voZ�l>��^3�?�W��c�J�^$�D\[�{�ך��t���Ї��d��8m�ݳ�J�mn��1���%�����w|]y:EN��Hn�p�W�������4'��?rO��vCW��ݕ��E�8T���g����T�3����y5�?7�94��iݘ���L��*׮��x9x�ux��S�9��R��F��(����CD}
��2J(��*��,��Qq9�,���&�a��G�|*%N�+�P��s��;��EŗD��L�IW������"��o`�u��U��!p<�zn[
 ��
�~�I1�\*�?�f	��H�f-�`��ܞ\��i��T<>w����c~��hK�q(�Q�BS��_���5`��z�,��~�]`��%c�,M>��:lb�y�X!����V��@��r;�V3)� ��&����?�����ުM��� �5pRԡ �X|��B%�e6�]�d^�'9=�R7_ޜ��ѫ��y,�OY�\4]s*���] ���ksR:�k��e�b[v=7��)K�$)(؎,�;ׂ��+JA�P|wZcg/4b����T:?z��O;ֳ#̊N��S7{t�zrm��Ә1q��tu,a#��VPܑz���C>�zn��@���} Y��˛��f��R�J2�yֵzXc���7�
�c("�A��p������ƽ��<<4�LXq~5��j-� �g�)5�m��8���L��k�C��x5�K
�'�C� T�v�=c�^>�����=��`}=7�%�a-�#,��bR�epJ�%�^�-_K�����
'#�v�������_�Òk4Yб�t�ܒSCJ$!��u�mAA�������(��r/��k=EA,dWg+��Ȱ��8�wv��s��-�#�a��ypw��O�>}�74��$���5���j�!�Ҕ 7�'�����Z���w���l��t���������U�qQ97� O���(n���𶒢WP��{��"膔��9���8��5��y}~5�W�ihB%�����G4��@u�j�0���z�r_�lѫ+��ܗ"�����m�8�����<;^���E!~�f/���^�z5�:a�IA�����-\\�IH�X�{h�_���z�h����[a�PU!�|/�3[�̝��oN��27��c��qx}}����2�B�7%�ޞ؀�$�t,C����]��q��n�5Յ6�,��������F�2��ſ�^͢�`%�_�B�����),���L�S�~]N����(p�t�^l ��k�B�R]�9�Q�ڇ�kk�_����q��ރ���駰�D�ŏ�ɜ���C5����o@0�$����z�X�4����cn!��R�lrjj�R��E=�Sq�$g��\��5\�Ƴ���7$�~1I~'\k{#A�kA�?�z�9S���#{{��4��p�vYq�A�w�1dQ��oN~�����a���\�>K���+)�����F;�>ˏ�joX��A�T>F����ܙn����2sTP��)¥�7��x�Gd��'){{�qb5���DD+��s�g3ܩ�\�j4�����~�삷���VZV步����_��]�����Є�C�3�J:�ZXוb/�'�B�i��t�ae�]w��l,�? �԰��J���4�Hl����[?�%.P�uy��G����9�s����y��*�a��:��){{�I��{RF,]ȷ/`�Fս �oC7�B�{�X]�sR���m��nt���Q(.QI�*+��g�]�nW��_�kء����50�����B\����7@�:���U'��1/��Ć4U�p'	`'{��f�,
pw}�p"T��[W�Ռ�_��
e�u��dv��\�.,�q�R\��u�j
'��!�:�R�4Z�ȁd��xp�I���p�s��咏�[���^��C�+����Ce�U��/E5��۟�B%�q���i�_*Ƌ�`�2�������#�T��Ri8"g=�ק{��FjO]k���J�{�-�o
�YY�)Ӻ�M���!���uh	�Yw�w�R�
�%ǋ���z��0���$B�V�{��������P�I��
������3C#��(J4�L �~��E��S\l'��t5E���݃a���p��h.Lu����M����P�7�^uDI��؟�Ǩ�� ]��l�6��.,l*���<�R[��*Q��FC�����=�"��m�;�.�#x ���P� s�۫�~U/��d�sZ�@�9b������Ъ\Be!�/�E�j��@F�Y
bG�G U���6�Oſ�Z�z#�я�La��S���e5���Ԓ��!?x��g���-�1��9�dhC��9�G(˥[6WS�<<�PO�ԲC�P�_�Ws<�G���/������D$B	Ov
YK�Ȟ��eߗ�����IO��I�o)����!4c�:�|�{���������>���y�׹���w��[����������;A��$h�B4����tsB�߲�̧�gZ]�h��������<��d)���Mh����;� ��k�>�����L����oϛ�m@�Ʈ��À5 F ���Է���S�4oR��D�����s�����&3?_�~�<i�Zd�d����&�%�E�b�n���2iD޷x��. ���k��q���۷N��%��ѭ��ss̓�z��Ɓ��<��,�v����o�k��5�ZPj+�IZ�r%�����ٿ���n(<r���G0���B$����x�ld���4�r��%�����������Y-����m��M@#�m}}�g��G��bmu���Z(({������k0_�HCn���C�g�5�&�>qk�S�����vv�2��\wr����ٜ�2��uX^��]����U�����x�����j���	h	��__��?;�I2ˈ�ό虔h���A/�n�ĭ�'�mssA��,B��G����x�m��E� 3x'w��D�5��וLb���`��c�D��� �;
��p�ϟĽ�k�]s͗#@����{�qS�G>�~f�σ�"�3a��io؁R4n�3q�x��N ���O�{������iw��s���t�͟S�t������rD��ȱ錄�����Ԍ,�W?��Z2� 朏8>1��۬���r�_��>V�k�3d*�k�'��߶m�)7�e���%���#�Ǻ>Ǟ�y����I���'��tR���	ٔ��R3����B3v�Ԝ $Q�	NNW�У���[�-/-5S��U�6��)s������תƺ6h�Q"hɺ	�6����Fo�\����	�5�:Oh�04R��8⬉3)߷>�D��\��c��)0���W�-�>8�zY{���Ұ|=ߺ�����_��V�=�����Z��UHA2�q̀���(��3�v�'o���6�=�R�V�d����Fp�eGh�F0b����%j~ V�B9��{^�@�*��"�vj��K�G}V��Au�(m��G5.��}���/��!#��.Tj�P�EeJ
�KG�<ƯDd�G�]Cb\7 ֕�,JHX�K`����9ڈ|C{����ÐO�;Mc�'Ҷ����\��i+ȣ���q�Abx>-b�Ǘ�d�70#C�`��	Bs[�O�yxd$0�41����F�/�4���n-��]A�	��X�WD�,�� {<�9�FH��.��-d�<��H�i| �s܁&tS^�&���H��cQ�	�?(�	��RoT�</W�XJc�"���M�H��&��Pu�;����WA5��	��oej3P�E&�^��0{�[�U�N�K�'a��nGD� �% <I���?��_b��p2jl��^/��K����sZڑ;��I@_o����x1�h�ޞ��FO0Ϫ��--�o'�
�����'�+D�pqb�Т�..
4�
��MH�T0�V�^�K��?KK��*���lM��,�%�`b%�=���ڍZ5(7���m�О9��P�ƍv�#f!������g���N���%���l���p���FM��0��>� ����o�t`�y�߫{�>��*{��m��@��� `�U"�{D����-<��n���3�Zg�h��8��f��J7p���<�n��Jɛ7���-�@����_�M��-P���px�����#	�@�d��11-��G@��|��Ex5���@+Aˡ{i�0����(�8F̗����˜kk����2ww�\��	5Dہ���������%�f�`�� �jڠ��ۢ��F_tzz�2�a�:�C-Ƌ��O�>]�f7��?Uu�_.4��d��E�Z�SPY`�N�^��I��Y��
�����Wϭ�[]�Ե��!�D�S~��e��֕��&/��T�P7�U���t7�+�ra���P��4�5�8O�u��hnֽ&��\p��>��76���y3[��||����n9SN�����✮� �������s"���X
PZ�e�0�o >�3�^UWU���%ޑ��\V�)�6�t�UNx��QPd)=c����~��k#���}��p���o��_��<x7$+�$�m߇��x��Xҡ��ru�f���H�oB����˪�+A�=�ba������P��	�$���9W-> ?��2=�`4���>5�HEZ�������W�LY�+��j~�RX}z�b�X�F	��0-��L�d�HIPQ	:/�&w39�\���q��wL�@�hyʌ@Ӭ�V�I)u�ַ��(� �����U2��fܖ.yg[�7�8�̸Z�r`I��xUU^To�铓z6	��##��3wuL���a7���Р(4�G��Z3�J���b>����c�nqC�P/�Ƅ"3��*�b(��6X���D��ꅃ��JΊ��d^�e�U[�6�L�l$c�L�w��b���i�T���������xU����C�UU��Y8�%�[�x9+骫�+g������H
����x��*e2�`c] 7a��gh�n?'��]�>��ы �A]1r��s�#������ã�%c�e���L�]�\�k��	�A\_W�-� 9��`e�{6�,���ήO-;5$Ԝ�b��j���:}��3�?�6pE*��c�%hȤq��t@d�"}[��8���=�6�w���a%�s�������{^y�ME��G$IV�63���X�����]�Lrs��IB�≸���g�4�]�W9969`0/Y};؋���\i�%�QA
�����p�dL�ߧܼ�,���Y�Ò~��x^E}����������DW
#EO'�����<-���>1����w�I�j36X3Q)C�rӁ<]����1�}�v.U�L���J���DO��oo���
��(�W��"$f�	Wu�z�uH�1 /3�r��� �@[Q�l?�����I/�[ f�c�>�d�Z�����mb h-}�g�P��`�&�H��EZil�\�A$�hvY�3�<�t�b�}����A;�Ryv���ev�ç�����C���.�F�T�)�9%�=���N\��8��W��:C��Dw��tv����_��(�]v�V�
5.�p�+���r9V;�����:�} �OI���W!ݝ{o��f�����5���B�8��@�ي���遣|Y���J���qA,6�6j��틛��OA�$��j_p|$Ş�,���F����r����j�X�|��K|�S�,�6����w�M�����R��>�� ��w5��*!�!N���M=���l��|p����+���􆧾�E��,Y�@�����YBi]�3QI����~9�G2g�`�4ꕠt�@�KDu��\��������h��$2U\@��c���CH0��E��3�#"r�@j<�!3_Y��q{&��]��"�g���"�б�a�\���$)�	��e'����I��J��~{==ZU`N5+4t�K���_�� 9�Ԟd�~����	��"u]Z��& ���ڔ�j���I�$�1����EP�m��c�Յ�:��-; R�V��K^��t*gln��}��>�Xv�x�����_�b�AV���������N������u��fK��>��ur�EA���&葠(�q���ҋqzVm'��!i�i5A+��;8�N�W�g��ۯA!7���sx�O�>Z�:��Hۡy���q�_���u��{Ig ןIT�}H��qA�?b<E��P����U�~&������gh��9����2O�xA`t�i��=�t.�An2Uu�5�t���:�R==��} r���P��"�b����H'N��Z��4BF��̋]��K��C�f"(B(���%5�ײ����2l~�~�u�L����ϻ����-��B5�m@����������J��ttQ�8v�!aq��
��Р����s�)���t�v|�/�Iz�%�!��.a�W�gJ��:�t ����N�T�J�(XY�83��I�wM�[3���9<�xI��\�)�x@jv$�����=C�k!-ш]�6;�?�(�oh���\O��Q�ǎ��lsS��?��A%�Y�z�
 hј�Ls�)$!� ��M����mon��1^6��,�Bv�|����/���q�(������ɿ��+�I}Bx��۬uH .�D?,��#4Ck 6Ed��x�G�:/��$=&���cQ���jS�R��j��]�b� �.]���(@�뢥.]�[{�6S8&��˽n�p�#�h���R2org'�����G}�m��6Ӗ���*\����?3S�<�� �91����܅��j	��E"	���ym�����=bm��+����V�L�}�*����R

rmU<��\|p�Z����"ĺ��'�1�`�*Xҡ4��i���VQ,}-���fހE�c�c����iy@�L�oԈ���̂�D	�d�Ds����P�}!x#�+�?pn���~�\��ut/�h�ǾM��/"�� ���5�e�v��t!G�@���^B�+����.�@\a�����>�MԐ�qCC���OU&�3Yh1Ȍ�?1�sمf�p<�_�x���D��!Ŭ+q i��]�m�'W�鍘!�?�Ek6�MAT���~�8���~��A��ö��np(Aզ�?778VE��7����f�DCf�ۘ�i�2_�%c0q�R�Ǳ-�lN�<A�8A�0󢢢��� u�'���u�s�<Y��B⨈ӄ)�I[ZM�����>�숑K�d�=�,�;4_��F ?���L�9����[���=TG�6e+�@����WS�It6�����Az�\:�^��Q��Y�ʀ��>i;:Un���:r�у*+!�S����(�|HE����
�+�������������H/��pq���ez����(� fm.�������~U�̌��e��A�6c����$�}�{����r5��}���ˊ���t�>%W�����@p+7��Ƭp�밑Y�^��$�=Ӂ�)��� �3��{����v�b��FD�SdD���;/
y���<
7�����~H��T�B������T����{kOD t�~p�A����Ac;t�쟓{�뚗��I�Vk��E�*�"+�g{y��1uS%��Ǆ� �@�= ��Vh�>�����!��|�q�f�1i7,�t�.gi1�����3j�x����;�O�;=�{kޞe	���*y��M_}��(^���.�*7*�F���a�3H��q�(7P�5rD�/�n뾊Q�����ҭ���,]e��#8�ə����R�{F���V̯��׍@�!Z�_v�2p�=��0�+bϵ���P�V�P���S$���'а�Z�pe�g|�Mm>_�Y�!jHN��`2Y�/E��~�SRO^���>��
לMm�Z�I|a�-j������n�2��݃�Au/�؇	��j� v�Ji����QM�G���q�����F�T'TF�����w����}��xDO~ϫ?Ad|���jD]@�l���ܯ��,i�F�`�a(�-�F����G�gi�uKs�� g<s:�χz���M�T ʆBc����ڙV������2+��X�:������2�`���4���B̤�5������}[�=��M��$���4�(�(��Ie�D�HȆ`�nƹ��[6��b���Y�t䚂O}�?AAr�C9}���<r�N{�^�KT��4�d��u�&�Q+�'�n�+mq���TF>��N2l׬b$9��E�1�~W�l�ڭ%���^M~�:��	U�P�������@|�^�z�*��&���tv83M�+u֯�~F8��k
j�g��RV/���xس����ՖP���)M�g����_&u��u6}֢�@c��0P�c��d!1��>7K�<cJ�*��?=6�Ԃ�M��w�D1t~����".+{;1�@G"> Vn��&4���%�(�!�!�i��=�	{�a�6�y���p�J�肐��>��q���f�����X�+z�Lm�+��(�,���v��5��x('!���quT�8����r���?-�&�����#��&�GԞ\�-qJ�<h�9E}� |T�S��è3|����]¸�t	����h�~�j"�-v^I��F�¬CX=z,��^a��-ѣ��eNG�&��p�n�()�iԈ��#�Ñ>Y����3	��ۛ���IK�嗇2�!����'nfiΩ셌T�%�'�P��.>mo^c��ߎ,�����o����Ȭ������ ��};�[莪*ī]{�rI�u� �����}i��XH^$�*y���g����G��7ծ��j"ʞ�s;��zy��s�Trl�7MF��2�>*
�m�b%�u�T"���U�U��G�����3�� ��?f�]��*g��X+�,�*%���}^)���j�H�鞮�,�|6A��:fF�������|�KR߈cY�xDV\�?�P�A%�k�t$3c��2�އ:{�g;^�����⵷;-K9EC"�P��Q��-%��m
'<d�|G3'� -S�U���ڝ��Po�C���04f�'4�\��s���h�Q����Pm�a��`9�?.*���XW�N/�|(I�hKϵ()�B��Ó$�nT_��S^������Ae�����f���d^t�[��옝��ᜡA� v̬��������j�CL|'>%�ToiBz3U䏴����~�B�9'��ʝXy�p�B͎�O���}jQ��[�vLIQ�T�<�qz`��bZe1�h##�ݾT�L;��p5wrr�M�Ǜ��������$+'%ER_Ŧ>�՝-*������Jݵ+M�"dz!/�52��vWf���C{�C
�n��=�G~]�~��>�`W�T)HkU���o�5�wX�7��;�o!�#������u2����P����k��bRH'��f ��q�x��.���/�B�ն��WK�AnAi��/]�2�w��|�77G��
��'(�|�z�G��ج�k��76�s�{���l)��ɬ���hA�J��Nn#H�\�k����F�O\7��8d�L0s��$�*��� ��\f��^��?v¦2[-��(~�Og�)�tO������X�\�~�"�dD��&8����
P? ���b|�� ��=I֝V��y�l�v�3�鶷ہxq�BII_hp��JM�n��b%A����� ��I�x�	���2�K0�\�	�QTW�H�����\KUU�"V7n'mϭ�=7M���J�κ��e�QudTF��-�	%W��9�*(��֧�O���&1��f_	d��/���d��"��W���,;8��Û	�C�a	M�b3b�+8�$2�9��0�^��-W�
�	�s��t�́�\��#�^��Z
.�.Nc�An�A�L�g���,�n?�!�3�4��H���������Q�ǝ�D9�uKjk�]�M����+f0R���i�#��
H�SQ�~�uA��ghe�t
�3�j�s��g��Ig�l��S�:/T�tu��^sy#	5
3y�x�
q�ix3�ٌ�\IKgܹ�,��ʀ/(5n*���=����jo+���.
>S)l�`�)�WD��W����͜Ø�:C�W�#�M�W����rF�M�=}�ࡔ���-����[�Rf'�d%�$����M�F~[e
v���,~��#�y@NoU&7�J
�?Օ�>�9��䝮p;�y�k�I" R�ab��:E#C��}���q��
���!����ʻ�;��V��<h?ݍL���t8��:Dam jO�?��eekv�Q��å��yͲQ�}'�pJ�p����lX}������j쾿ˈ>:�h���"P�?t=Aj��p�[�]+3�k'�iWa��3<'��^̓?w�	����2 z4�K� 	#��sm��s�s�Z���nV=:�?L6�ܹK�3�l��'(����m�G^�$����C9NLЂ�]�yx����|��+�Ꙥ����{�٤O�:ҧ����U˻0�qf@n�$��OC���)�8(�O\`	��݂oF�V FI����P�㱁I����cGlA튔 (�b�E�p�8���Lyc��P�i[
yk_��$�@�ޤX�:����� �`�Z���J���.���:f&��?_��8�����W��g��b<=���Y�a_�djR�{㷪I4��abYC^�����;9�$£\�q*yok�6�r����_���ҷg]��5.���C���߃U�-�>�-m@��8�$:%��ep�!�*>3<�k_5�VB���C�J��|f��{⹫7$�v.�ٙ ���>��_~��#q���=H������,R����Y+��0�:c%%�kR���"��q&����R��V�ww]�5�K��,KD�LH�[切�e�{��&��`�ݣ5�G��|X
'P����Ư�{���@��Hd���C�R��l�HE��(�F����^��cs3��]�������E�]
Ww*�eS��r^�T������X��~��F(����>7�!���w�����Ak��O{���	����:jc9ˌ2��o��ǡU��O�9�c󺐡�k�	]���'�^^�3c��L}sL?����}v����ڙ�w��ׁ����B��<�����Vh�(�t#�	h�9�.���i���,mjT����������������e�0�����s�`^�6�u��k��.P&Z挄o(]��Xբ��h�:A��v#��v��k�h8�h��7a\y�g$!��Z~��6,R��3_N��;f;�XyGH%�
<����/��ݴ�)C�v��J3aJ�Lh�&�2�k}1SpvD�|>DJ߉X��P|���R��D��V�F���%��	ʨ�A�Y��{H::Yr��L�=��[/9�iv�ۛ0������yr���ӏd� ���K�
8: �(�.�D���z�#�J��@膦�v��}v�=9�����9�"-P�E%������<��V�$�;��ߍ -y@�.�d���XHXH������ѥ/cv����_�h_F,�B(I���Î�Z�I��,~�u�#'p�kХ�����$&�,G���cT��GB�3Kmnp�z:���<7���_]��&��'T(^M�/��k����#����u*�9�PE�����GI�F��`gCCA�ngZ� ���S?j�|��Q�K�.�Qv���g���[�g��Fu5_c걫�t""b�\Ei�:�t�킵�g9����ܐ�[t�8��}��U�>���RR�w�JO��9�x��.�EV��l�xR��m0�a��9ӵ��.z�N)@�w�cJ3���eR��<+l�:�Y�z�2�]�l)Л?�u8>��.#��g���zU3��>�MQ3r�nRi� I��W&�RgHڴf�J�� Z�������OW��Y�H
�����^���?U�	rz�U�Mq4�^M ���l>A����֛ޙv�����O��X-*���kY���Ŗ&uz��6�yA{�)wj�O3�k�!�ÍTң�>��� ����X��םi˰њ��K��Y'zJ��%� ~����o�ƛs�������r�~��t������ � �Ł���/(T\TB ��iuY�۳�����$1΁�_�F���B���L���JU�����	pHx�ZM�޽Xn�<���^��m��4�7i�/k°�� IR�1f�Y��0�?AE���������~���7fU��ɳ�-W9��7=�Q6���8	F�;��xڤ_L���&��`J��������ԓ�F_��Mv���F�S[�U��bi�T�E��0��h�A�aYQOd���@(���H+���Gg��2��5��uYY��,��˃ڒ�dj戴���b��\^�ܽN�����+?��Qk��F&ޓ�\�ذ}��"��an����(�:�O���������/xZC@"�t'V7�NqEE<-�E��O�hu^���ִ��%�z����:�]���󾑹ц�s�r�d��q7�w�DYAO��Y*~��͑l����D6D��5�՟q��M��y�p'�?�2$g�-.贅�(��=��Ͼ�z�	ݹn% 
D�g��]�����T��`�yR��R:��n�m}�_��@��!�B��Y�d��O�����L }�U%��i�)<�a�e��P��l�IՆ~��ڪH�cý�ӳ��js���H���uW���J�s�fSih�����d�'�'V�6�O:=�sѴ��Vn�gOH���S.]Q���ŵc"��\E2�!���P�D
1>T��J�	�7\QQ�tGyz�h�ط�x���IHx����D��<�8�Y;.���m��jY���o�[���Th�NF"��cSg��5� usS�ڛ:&th�cLG����$�-$ޅ��n)fҾ�1�}W�nx���u��oa3�����&Jؼ����qz���q���q��3kNNN�T���pu�ίB�>�'�$��t�zh�G���R�:�X� ����Zm�ԝI�ߢ��t�9�87����m-��CC�=Q��' �W�<c�8v�wC�-����C��]i=�!+{�E���G��PgC"���Y9k����ኃ����[1��Wĺw�����5`���Au+�����@o��UU�ɛ�roS]gZ3��(�p%:'^(yCG2;A�kT�W]���1���v��g"�ZZ��M��4G���u���O����gĭ��Bѥ�{�p����|T닢�4�'����i6�a:El�N6Vإ�~4�/b�\��}*(��朚��r�'���^�}T:;m���u�Y'�dF���Շ�A�K�k�%1zz���:����B�H�6	j�.u�8�g�/B6���<�_�	Ci�]�	yVp5y	1��$_V6Ԫ����.#-�{�r����p����b��*�7޳�)f��[������.Ǫ�t ����vA�Y=0y/OZ��YR�/q�M�u��;�ݧ�ٴ�#=c� �
(�Z�d*w���"�6}��Ɔ8���y�V���B�f]��S�jlj7J��!�c��kލ�b-B1=��(��@�t��p���n�R�´�9)Պ�����K�V������!���̀5ǰ�m�i�g7D\"���L���{��B�-����[^�����ٕ%B.�xS	�fݚg�;/K��K��6��&ZZ��A�2����&I��c�6ixkP��z��MW��2<D�E����r?���e2gj���� sQ��`J?��	�������==��G�a�'�d�1
����g�	���XHz���,�6��!LK��{��=&��3�{g~]��n���ր��޹��_��"w���hWE\��V����o�:�Zh������l8|��@
�J��P�	$�S����p�TTe.�.s�34;�Q}����-%"�����K���XB���fF���V�a5���r�lN}]4�R��5��gE�!�'�%C/͌:&g��_��x�{B�DE��5<eWh�$�-�6%��u'��V�E˝�i�ˎ_���W�j�3]K0s����D-o{��'�bz�>�N�@j\��ZB&J'��D���g�G�~���FY8j�<�)ФT�`+j�R��"ٝ9�����Ǧ=��[I6{3��;������I�l���Xj9ȝ s���ތf4�T>���?���c��I��^x�|��q:�
���� (	�W&l@3������h�,���mE��Le��K<�!?wN JL�@����t�Zg+���'p �*4c�<��-c>��O��"�[<�9��%`��h��Vn4�0Q=A�Y2����$�-_W:X���յ�{\4K���/֨.�M9$�g�G�gK�a��I���<4j{�m���a&�l�����C���p���~]q����|;i��ى&ݹ�\�i��M#�x�����~t*~<aI�B�s��5K��A���o<�%LL��%�����W�4�wD����E5��)Y�i�j��������vHl�>f��=��b\G�<�Q�e`�Emy�r{{��@妫W��G�G���"�@G�:��h�Y�"�&F�Cw�fI˥�վ��c�؃�
�;���Ƥ��M�����u�%�nyU�YA'X¦_R=�Q�E˩[5��g�b��5[�[�F?�h���=�X6�y7SR�;���I"�M����7�Ӎ����M'�xjgO,r.��s_�[cS�z݊�c�������E>V_��X����`Ե"w��c@=�loV���Pxv�خ�Ţ��-�n���	���^V���/�䓿ہ}�󳵍XD��T��ms��2�n���
���✖�If��uta��^f����`��?�^xTq����y2ZT�ΰ@��qѕ^����/�E��]�g�,�3�Y�vCٮ�Y���t�=�y�Y�qt�Iٯ�g'��&��9o����l��_T��)V�RhJ��4���n���H�L-�G)27s�ǳ:I��Y��I5?�YR�X�F��\v���;�S�m���k˽�����;9�C���7i�]���8歕)�w
	����]u�V5z��`���	BB��}j��Rô��+f�~@j���a�0�!�N�g�4Zv̤
�B1]���$,���f�����e����ە��XD@��]?�e����綪H���3x���q�/�.��)_m����͎-��yx���,�(��1s�Ǎ:+�C���K�O�Z�W$�F�*/�y�.�b�)Ø�2��f����Sa:����F?���q�G~��D��9>�t�M4�v���{���#r�	�U똩�c�ʫht�g�u1�x/����es�h4��L�?T�{tnt���v��W�%Q,��vo�N/Ifv���{f��;L��fVE���G�/��#�.����"�[b��'Zj��?R�\��_�c���U�* yKmj�|^h���L���U��I�&P��̊�}�7z!)i����Ì(���s�Z�z���7��uUڽ�o�3+ҿ�&�o��j�|×��b����V�u��#�������&D��nX���(����_�����v��jm/����LN�n�m[p�bnqzǏca�! ޅ鑹��%���������h�5��E�������$�Zw�Cَ�/�uh�qU����w�2�p�Xտ�����k�Ӳ>���3ή�t��IО����W�wwcS�,ރa`��dㅫ�j8������[˅�鞆0�R2r���Jע�x� ���x���s�+|�����a
�M��/�.z�ݢr�G�
:ť_Z��jǡ�eǼD���%k�WR�XL��f���)��e?��v�aXN�mM����-4'gM�L.���f���m�4"x�z������
�g<���vy.��E&v���{�X�o�"�
���0�SJ�]f�:3�8�[��%�6k&�9�Qa�|��kc�VK%�� M�_�0�y-7��CW�Y��)�M��w�����#*X)1���x(t�dЈlʉ�~��]���)y���Һ�3���wʷA���v��=g��[A���abڌL�F-k:��-~�Vqyy�9V05�Z>�:l�oG��Ȯ�f��h�O��=�n��S��R\���?e�;n�&>K���v��(�`IE���_���i�=��'*j��9��d�p�
��Y��.�ԯ��+�Soe�)�S����.A�>�:�p�Z�����5웳�ޡ"���έ�'-��蕷�rI U�O�{�*�������e�������+����\�v5Z[Ӟ=�My+�E�se����4ߵ$�?eEభ�1��
KI6��;C�睎��YF�=ȜBjZ�� ���~��
 �Ȫ��#̱�/�E��r8k��`G$Ѵ^(���:���TI0���F$�pa��b��]&GDd�$�x�����<�OMnw���{�^���z�sjΟ58y39�>�!22s����W`�+��b)��v?����X�a������e�������|�zVs��A���!�s�o��v\L�g�	������2 �,ƃ�l���š�����;��	����t���۞c��7Y� 'v��ΕK�R�7Qҷ�w��Z�I�<O�mɰT�M={WW��Ee��a�[�K_��b�>��y��DAH�<e��y�:�&=#��K�2��OJ��s>M�ϙ�.�x���9��P���s�#�; q�1,����KP���㷦إ�,�Ym� ��+ ����M`*6}N����԰{N�[2��;¹jtQ�f�-����}�B�[2F��V�h���2At���gl��;׍~m�Yu�+�2�	���K!W`H�[_6��EVk�Yb!���D������g��;�[��.����q9�n���(�H����B��A^�����I��=l/�D��^��h�cQM(�_ZcbQ�;���CٌOm׻�5N�'J�lm#��]�B��f	������4�`"@�#��o��8j����}�x������Y�W����,y���|�66��J{h��Y$���$�����5�� i���G�e�J�}�l�uk�4W̻�~����O�.�	�n��Aײ���F5[�z~�wo���+"8,t��e�7�_��)������}4�1�ކ�F�A<pP�,.?G�ï��?�8$z0��,u|{�|¾m�OR�^�pFb��(�G���<LM�.������L@� ��?^|d]����n�Կ�����J��1�(��B�o���QN��f����e��T���h�ҳ��E�]�0FP��Da��i	V-J��u�»�k��P�ɛcyN�Yx<Sb2�K@Y�M:�w�n�"!sse?z���l��L�0#�'��n`�� ��G�&����<�������߶&���4�h�<�̊�m��20T95��i��?OH�	�'������}C� ��h�'�s-(��p9(��gM�_@��30N2��͗F?�65GȮ�,��r��3Nb�(�V��7Zs���*�Q�U�F���ICޛs�����c*E�d�$iD�f�A��߭k��N`Ys�X��
�r(`�H)�F��Z�Z������X^^ŝ�&W�sa]Ե�p��T`�I��f�+��v6/��aR���O;bG�%�h�����`K��X��d���h?u�|���4�"�u��+yC�س,��Mx��o̝�}�Ǖ����&�0�)�$���^�ɳv�u�K���.M�D���5}�������gM���[+$��v[/���"�I��h��w]�}g���N]�w2$��@�Zu��P.:�wf3��b}@������D1	���k(QS��s{uOx���p��Դ>{�ë�n\.�����#�"3�#,Z|�i@���x`m�LJ�M�B����kتӳs���m��0X�A��l@0�aD�Į�0�~��0�[��7����Á�2S�i�&:�vmo�i�?3��(��ϹAf]��B�|��-=�dc,�� G��+�*���TJ�53M��Z�9�&B�V'�r$<��ڐo��JRe���M�F���E?O��/fћ!5��fW�������9nP*e�U��"����6;��Ђ�2U`V�Z{�i ��4��g��У�/^� �� �{J��M�y8���^��͗;�B�L��}P�5ڊ�� Ņ.�e�T�2�5ຜ��YJ� 9l��L�de=h�]�����rt��g(4�@���.���4|��ϻb
�ax !�Y]����T؞)K������K_�g6�^�G����4W�6����wA�(��#�)[���g������z�a�M���U�*ӵ�?���Q�AP��|��|�P,�m�s�Ű���'�Vj�l4� �x懟T,#��+F��L��O����^�!1,������ɲ9"Iw�O�����9����Ui��t��@���m���S��k:sOTc7*8��}��v���u�����zi����Q"o9�=4>T蕬b{V���?�ԠP�����q�O��\n2��?w��f���+�-�=����p׭ �~���
/�k��A��ݱ���2�r�ǟp^ԨK{�Sô��8�
D��fX>x�>;{��0b�r2ܡ��`\���5I+莾��������֟4=���L�E[�E'w?�V/�"}�$H�V�؊�O���l~.�a��2VӍ�s����ኗ
E KG�v݆Fge!�n̿,d�,�y��o���ꑋY��k�]S��8����&�xg�W��WCG�v�42�Z��SC�����	
ڱ�d��u�uiN^�]��L�)������ኙ1̠��u�- ��9����,̸M��bb���ݭ��[�ڹ�p�^���������rٿ"JO?�^u�!����|��G�;���.~.7�r��OR�X.*���c[��*�	���?�,�M���wB�g5���Tf���z���sv�����Vπ���H����_����.�gF\f2�.�0pz˨.�|� �z�^:f��Z (��i�E�j����!G-3x��c��9Q[���kz�<�9�Ӿ�З����,'�Gtq=J�S��c|]�����Y ���;��?|�����$��p�cL�ԅ}8Y����I�B�^@S�:(ߥ��E �k��$�۽�{�E>����B��\P��ڑ�D���g�	踄X��%�!�h�2+� ��%��s�� �X�4��ZaUl {ST�,��C����br%[��z�nG�O �[Ԧj�.<B%:�����%�t�ѭ�5K��Ǘ<3�К���,����fE�ui�����"..<9e��[c�4��u^;�ȅ�+{�[7�KH>�QLt�l��lV�+�@/@����+�F�JA����9P��Ũ�֢9�k��d�(����)��i�G�� ��G�9`�Wt~�͓Z�E���H�\��!����~�Y��*�`$���ʡLY��2��[3�u�X�,П+B&<�VG�����O�s�?�����z��1��۳g�f����wb}G�eM���kқy^X�>��Ӣf��(�\{�sy,��6vT+���v?��*)�,?W�h�^�8ُ���$ ��o��-6�2�g��%*�jo��63;Vcv�����w#h),���ؗN��Ɖ���������`�{�9��2�
������OW6H�;N�\ u�tZ�Y������)��j�%��D��u��7,�_S[@ݪ9�`�.g=��=�H��U��k��B�/̊�K���"!���@�M�� �ޛE��-�ܭvl��Z_\HcP Q��R���~�S�-�r�_��Ujm=�.n�/��'����#т��/���������nra�=��z����b�h�@7��ܕG�.Ztb.lV�\��J����܎��~$�l�b�yV�ʎ�Zb:<��~��z!���K���B��y��	��7m:Xس>Oڒw+�ж��J��w��C��E	[SS:�<T-�U�����a��>�X�G�v
�h1�����쇊�"�!k�N�g��N�>RYX�'�W���|;��`>fӯ�p�W!��R��r3���$_��Ix*�X�ey���㉢xV�ݝ��%RO�~��"�&�w��<��gV��=�D��W�/R�:��������vB�|��3���~Pn휋/�a�g�O�a�LN���m�F�)��`Y*�R�ߝ�0�:���{��#��d:*,I���_�uP�n�'�}��f��Cy���+��no+~�'r�z���1ܫ�|$q5�$D}�U���)]��;���:!H��?�^7:e�tV�9�ś&>�$�\��&�2u�4	�R���K����v�7~�ڐ�����6~o�����$�Fp�aU�q���V�i{��;S������*���!u{��[��s;��j�c�d	��f��V�&[5���:� -���ocF��,��
�����}4�K�(X�f���-(�����W��V����57+|��~�U�|3�(��q3F�Ĵ���m[�G�0A�æ�x�����p��rč��;��_:3��t��p_�tj��?�x�+1i�7G��ޔ(��եy՘��?T��#��,i���l�!A#������8��B�o���?Җ_y���X�U�����p}�?��:,��{DAE�E@�AJRQ��.II��4�G�����Jb���$�`�y��<����xyy1g���}��^k�9@�}y7;Q4%��3�\d��{��_N�^���H�B���}YeX���A[�]峐'�|�`�Q�t� ~Om��.wP~���?��אv�T� ��;dږ,rDe���>�CN�A+?�y���si�,��%��n{<�9����%� �z��|�]s4�����ǝE>��a'4�w����@�b����H/�X����w�		��w��G��-�O�CK��9������8�8f��P��G͞���y��8�o����N\���C8!p)�XZ�f�r};��w�$������z�w�R�|�~����)Hv�����"��~[GGg8�pe�G�bz6h��_��q+�mY� �HA���?{�,
nE����;.�U�yrs��9D��U��>���T�Ĥ �,,��֨炵ۺU�}c��	��[<����FW;F��Eo��k�V�����՝��J���B �q��y�|�|S�D$ dθ��^���ɣFw�ݧ#�n�ē`�.����_ 	DO���K`�ɾQ�n�U��.$�|�:>B�d'bE�y��6���� ���m�W��v8���8/��D��]�`�Z�v�ی�:�f�?�6C��Z�YN�����
Џ�s0��s�Ah��}�� ʅ�ȩڋx2�4���홓x���ס"((�����Y����KST���(�� ���)������$��'�}�-�j爇�W�8pؗ�q��FvM�ģ, +�?�"�Lz{����%�漨�]���!Ga���^�D	�WeO��Ou{a��"���*��98t��!HV�exwP�k1�޿�y�~�N��YKE�D�����{b����E0C��r.wb�;�_�z=��o+�����J D�����R��r�
ѯ�Kɔ���,Ѐ�M�,��Fx5d�O��ѯ�zH��������l����R|<�V��+x�����Q�ӧ�������..[K���	��G�Y�@cQ7��2nm�+��ϧ���c��&v�:�����{��9.-�,SM����ҫW��h-�:�N�$;�3(k�������e��*�?�j��WZ7��(uHT�^��P����)�i������э�*=���K��/�rfڢ*���`uwO��)�7q�svW�'w�"'�9�DbwP��5Qk*���%*�$V��l��)f;��9{Jٳb��N�c&���,���I7�+��4s��p�b�cwm��E������)R�YςkJ��w���R�0��Ώֈ�xy]�C�@Z{ըw4n�7�����{����>���xS P8�}/"��wB6=ȇ�2�� )9��e:<����n�?C��\a�)w��� b�x��X���+���C��}��.����h����dw�;̡�F�����v��c��>��Κ�+��T��2�_5Y�:jE������Zj;�Alnr)�^x������[2{}r^e�[���1y��^�%�D#1��p���'�4��o��NI),�I����iHx�̸����6H���2�"���>���c��=S�����j��eW����e��0K.���"�:Wٓ�M���J,���1V�8�l��:�<4�@S`���s7���ZNlPKK��5�3;��!����g��ޗ_l-W�	��e�-�Dॖ�N6,��o|{���d�<�"���k��@r�����ƁCbخ��|�T1&��UN�7T%�Zak��VX�BBO�1��3�x��'����Y b\�@3�()鮑e�����N�Q��Z
��(��jCYWp�R�Oi�����;u�[�	[��$�K����$px:SH^��
U�Jt��{ �@2�Z�Y��3k�~JH��H�_h*#��xm��)���&�7���f����V$�U�
xl��y���WM��+=C��+�����ѸO��cw%��0GNw݀`�w|���|quS��`�'5�E���]vW��ĩ�	�K��̉IT���e��w,O`��,cG�����xKH;�x�W~]����P�}8����p����C�~o^�vnع���5
��2�Z�=ѵ��v����>��}v�1�L����q����sj�!.mΫM���/�S�J�����{U��0Z��g2ҙ�$jf%P/�%VP���O��8+��w��L�MX���8��w�A����aQ������5�C}�wJ����CTbי( �m�����Y�%��e��r���;��F3�$��EA�-�/�E7N@���&�]M(�C�E�"j�X�#��_Q�׆�x�"73Q>�%	���Z9�����sG���Y�1�9�wx�-���w<���-XOXVơa?�w�
1�e��+VA�49O{�#~�J�b�	��>�1��ןg*�������@��g]_�����L`��֔N���(�(�*�'�i<�3?�<�bp�EII��.>I��3���l5S��	œތQ���[fD}U�f��x/|Z�<ۢH�쇈�v�����\WU�2���qy'_Ֆ�Q�O#ݼTf�h;��a&A�x��Z�е�_�W<��h��]�7��&,�o�-�.��g]AA���ݼ��),�m��9c2�9������lP�f�I�y�w+�d�zr����0㗞������=�����Ft$��R�/�DC����Ą���7��jj;�����~g����xcj�7,��r>Np���9ahdc9 k���^xچb{n�c�O䔂N��	�p�ݨ�:bG�MA�bR&�B︗�[�5:�/�)�\�d*Y�'�{`�:F?8��S�P�e��V��V��\/�]#Ǣ�>����/���_��-�bf�����7�"R�I;]����Q
~c2��;���)�t��J�B��]bV��.�(|��<e��2fw�T8b/39� g�Aby��E�a�u\�2v9}8�8�����~��FY5�h�0�w Ȩ��+�A���51���J��ϓt�Z�;p�P_��b"��j���?�1���/��2����:9u����U�?]5��YTFu�mq���x�[��~^Z���X�����J�M�Z��]A��ԲL��5F4���Y��W5�!cq�,rq^�>�������3K�A�χ�jČO�u�\f����t�ݘ�Z�����>���QSY��W���N��գ�Cp!���dC��� *M
�X�P���XeKdP?Z��1P��CQ\�zG�lN���
~�ʯ˧�&�-��=)�m��%� �An=��������˲�w8Me	�����Hs+�o�V��*´�486ۀ70v}��g;fџq�Ӱ����f�)Gwj�`�խz��8R�gh>}S�KC�g�</d�
;S�����䯏��e+��'"��R�����,�e�bK�v�-PU���:�I���V�i���i��n� ���J��K�}�����\O��9�Y�^8l=`|&���_%�]��j��v�\�o�s�F#&�����0�g��@�����}=��w`�R�S�p��� ����?b��Io�])���Z�N�׊���`���sr��}
'yg�;�ٸ�\ʅ�.�
{W�Ϫx�H��07�v��%G�w����]��@"�R���+6�S4���\�<X��<PռB��N�TV�Jp�$�$=�P_?�q�9mɷ�N��}�����q$`.����un�}UG$�sGSՠ7O��A$y+^�K���\�~�|K��_��9��>M�:{���͂Ad��M��2O����Y\�������5�$��АW�/K���w�J��3��{�l��*4A{�|����^fS\��ɳuȬD��&���0��^����Y���M�	�Zf�������,g
Ҹid�;u,��'M~�p\a���D��v�!��k�X�9j'����D||Ӎ��x���Sq\�1G4�尠�Gʘq�mX�q�Cx�+�s֨�^lR�<3��Ь�<Eqݝ���҆�~U
g��]k$+�#p�o��=ӼW�&�R5va�!/򉰌C&�↯������B�~�ă��;�`0����GyEu�
��6�`Wt�2���Ts�6�v'��=����ә@�"c�w��쌺Ys*%�)A�L���!�7�0b�z��-�-2x���W���Xe�0ԉ�Ɉc�}��z?���G}w%%
{��/R�A��9� %:��j�����M��g��Q\)R�Mb�ų�]�aY�qT!��Ƅ�2<"W
q����%�WM����8��j�8��UvÛ�DA���*/���	�XA�홣h�z��Ԟ5n����ƔI��ry��<�i .μ�|���}֫0 ��I(���!b�<s����J��`���(�ӿ>U}a<j+1�s$$��#��Ӻ,4��߅}�[аע}��f�`��s}�6��;��M�3��$<�Б >�OQ_�y�Zԏl{��{�z�����
��9}9v��%+M$���p���E/����N��N��kL�C��H�Гn<cX�\���/�L�����O�Y8�pA�X�wp��~H-���\����pض,q�/'A�:�����V��5��:O�u�vG��8b�綦6{����R���w5I��<����l�j�ɧg�R��P~8����V����/e��t���w3p5u�@�g�ӡ�9�@,{��>.�I�����;{����"�Z�?��/s��@('���K�h �8w�K��)�-�`�uw8���"^	e[%~�W���q�(��\i�	�J�L}O�34�oPk{�;oࢴ��zN���We-����Т��S���%�¡�{)΅�ӧ�45�֩�҇�@��'�����]0�{-f}���>�:��}y��5i3�<O����a���rx:0���w׏��D���I��<�o��-��ځ*�lo��0����� ijz}��(�R�ng��d����$f�(���浑gf���;ļ��	+1�_=X��8Jb~���/Sf+Z��-z%�(�~,��ܓ�n��V��y��N�:�"���K����vW�C86#ޜ�a����`d��f�o̵��X34�g�JM��<�=1:��<��'"��jC��.����6�;[kyu���A5T�&�f��3K�$�:�<���~ؓ�a����F0�v�����)��~K�SV]k��@��s�: �'��qB�L��R�)�eII���נ�vKbȏ3!Rqhqw��sU��^����ZyI�\�k��,w���s}�v��5^ޛ+�Z}��q$
l�FL�U������
�sP�5w� �@ �fd��Uc��0O�/���Yh`�1����b'�n���=Ą�_2ߎ.�ogbFy���k��k����F�p+U��qy��m��m5v�=[S.U�%w���g�4��㋪v�P���}V����A��l��y��q|�}� �~����)fq�&)��?bbV��H�)*�v�	$Qp�yRC�k>,��q�ȴ�CnH�t�D�袡-�ӫ�Wi=�3U��$<}�'�J7dO��s:����T��j��� ����>81+����i��S\O6�;�BBE���3��g�C��ߒ����։<�{M%���*�@���O�6�E��|�Xp�z�i��4��x^��T���43ZZs1�}lD�>�K��~#��)�%v)�W�j�㇘`�
�TX���1�c����G���}wR��wܷ���ǄF�ϷX����r	l�8Ծ���78`�A�柚�i\�,wAW�vKH��M���͐��B}�.v�c�ԙ��7�+_����s��@�=	n=�d ����.y�V$�ׯ:�S�L���=6�N+Z�A�󘔔%���%[ِ��ND�,�(��f^���bgC�}|��W�<<$@>>�sU�Z�A�z���F��c-9�9d��m~g�^������Ξ���e6�s��}��0��EF�Y%�a*�� Y̛�{�rE-sn�{J+EI���k�AH��&�F(8�Dr�I�YX��ry��h_��k|5�ס����ָv�_��9̲̔?ix��]w��Ꮾ��K�^�A�ё�l���b�ui�'}�c�ʲ�������,y��A��������w`\�<`ld�G���NJA���7B�5^����Cc��([�޷�458}����:)-k��`��qGb]8�ɻ�2�6�5��
u��]�|�-T9M�w�m����^mT�ij�L.w��W}=��(3�@�X&k�hZ�Ϳk�og��4))(�(>`�&�z��Vj>C�x��~؛�5�a��\�d=/
2=�ʳ��ۆu9gS��\��R�z<�3ē0:{K����R��X�e�$
��>��Ii��b��X�_�0���Jӛ��{25##ug��4=�?:�XgG|�Av�kp�Khjn)�/�/������D��*Z��F��H3+��6�^��]�ޢ��%{u�%�l�%myM��c��K�h����w�C�����^�m��r�I|q��f�7�
�r�~F���;wB)|6z��-`KfS��õ��ʒy�n+s�����.^QZd��춓E�Y��WT��G�h��r\z��h�_1
@A-��އSW�\/ }������	2_�e�Tfi����n2���v�b)�Îu;u��.����r��v���Aibۻ�=�t�}�P���ۯU�K'�|m�)�:n�q�ʬi��Q�P3��R�I�7o����E��a��-���2VG�������q�)3��$��F�b���J��5̐��UTvTV8�Ȟ�:8���П��7��=�|�C�տK�,���X�k%��5�X\Y�y��;uqN۞��Sx&�+p��o��Lo�0lMLJ�` �ԘvǑ����`H�_�ў�f(ΰ���#��x�ksV>$d�ͽ㞰��JQV��#Z6�C_T_�|�  �T:H'mpl�m�]��u���Qѕ���C=�g�6����}�3i߻Uֽ� ��^�w�d��B����$��x\^���v4��26��_;qfk1��ˇ�7��W��t���,�gZ���ΕTf$�r�V8�ĔHoo@�/�-]�FS$1���#��.�a�/N-t���ר�_gnn����`1�{XB�{�H��cԡɤ6��
z�e`Э�bt���4|�#>��&��M��ZR���#�$5��Z���YB���A���b�7d!��^P����pe�`��m`o���ߊ��;Il��N���Գ�����ڗ���öRQ
�^x*���fb=���Ԝd@JT��	��#A��c�as�X��QzWG��v%���z��d��U�ڟh�H�|��h�M:�L[V������_珗{�o}+���BL�YS�_�̙��.�F�!S����N\���@,FD��K��{e%�&+�be�q�[��2mS��Qx:�)��Y"�@�D��k���-[�|�"�C����4��C�AC�)�[��<Ej���������	�,22[n|�
���)��[*/ {��O��MA�pm�e-��q[b1w�z��P��k����!�y�^[JZ�&e�l84`$�@����|z�~N�IH���.�w:�Ƃ
�;��JA'��ꩃ\���)���"g��<�ge�x�&�ֽ��&�D&�./��o�6��E^������gM�8���hA*��Q���͑r.�G�6b*	�
�X�$b�RC�<��#��B�W�]��N .T����xM��fߦ�c��J�:V���:띞���M��(�$�m�C�^�{Bi�I���>��q���7oj��*�;�vwo��^�h���6���v�Pt:��x��1��W���AQ�b�@�[n�C�^M���Ҿjj�4��d����^u�6:�8�E4+�����N��Ó/G�1�gUC�bbp?�e8��R��~�J����#�T�sv���Af�Hsy�{�>��Z���������}���o�[O�{�Bng�@��ᔡ߅q����?ȉY�+��B{3�����7J2?ɚz�����M�>r���׫̭���U���RD��kl�˭��'�XU�UWΫv+x|~$)�VOl9��R��Sw[��]�S �Z��XϥãI��n���"�;�U�P{�
'' ��M$��7_`�(�Փ��M/�;3%�eq�c����}x��j�A��p��ҏ��X���م�R0����P��.y��w!ZL�\�9IM�#M٫�7y���\�����N��YZpK\�����4%Z��>"�DrI�|yW�� �i�a�ŶNV��;:���է�
�a8Vi'b�QY�^Y���(I���lLW�9z�X�Ծ��r�ۣ��3xѴBP���JK��+f���5]�c�v�ݑ�]���W�F����R�X�%�0"�M:)vv�����#"�6��*vm���N�����ط�x|x�>�W��싦����/���9�+�����g<e�8ȂG��,��	����X!l������� �e�ݜ.a��NQe��s�����6&e�u� ;����A�{>�� H�=�֧������K�A��-#b0\';}��g�8<������p�*�;��O_��kW�K� ���7=r}N�EM��51��L��NYD�<+�|�.� ��V�J���>��0�:���R��1��ۓle��X���hkda�b|T��[�Pw�M�?�������xqj� B�cH�/ՠR��ZsߌYR�g,�斖�������ɑ�#����J.��҅w��
�����֞nJW�u��\׽�(A���½pF=G$#��D�����.Wt)[�aW
w�~��(ߜx����{T_iڮT؎�_�y���J�F�����|C����Q+}��
�ز}v��<��[�KK1�4}rvI���cC{��O�dq�C�>�h������V�xEݘ�|������#���('�P%�`WEUo2�p��Q�䴍U�/N:Npb�@�
sԻʭ���4��	��&/ ������ߋ��������t7��$��(G���W7��yH��x#�q"pKe"�%��'j5_��ks�'���D<6	}L�:.`�GP��5��.JJy@C��ᖤ�O����� �<5#�ظ�k�Z��5��Z���2[���d�DWyW�U���;�;QR���x��^�`�(�l��^��d�ڟ%���Y�@��რ˴��@Ա�Y�ch�tJ�x�R�R7zrjs������u���K��q�N�\i۱nq�S�(a�d�i]���4��Cv�?ޮY��bd8�L
Q����Ȃ�Ȯ������_%�ϝ�/�Q�\f��{�
�U��՞*y��f��a�6�@F%������U�D1os�+���R��E=��{�G9���+�lA5�z�ѱ�D���)Xtl�+xCQ�h|؝̹>f�Ha�O`��(/��Zg�66GZ%�&���~��
M`
Bed�b����MΔ�a����`qA �g+*�-�ndx�_~�����.3e���;o�������k2����p�	��>�2P�9V)�����-	��O,������Sz��i}�P|���ze��[wY4��mg7�C(�J���{�3�- C(a@qʫg�����;���3�V�N�*����Z���_tn�^e��'��~�����@ӥ"����ROv���Mi�g��#�����
jNO�����l�����b���7" AB����m����P0�(1|ېK��Rc{���a?�kܙ��t�_7�_5.�'���"�1!>>Z�N��"����G���+�<�[v���
��.����ևd]����+���	�Y~Xz�F|��S�Y���;�k�]45�qC�O��a3Ϗxy����dd��t��Ź�����L������ԅ|Gu����B'6W��.��j���t��h�i��a�U�����r��McuMs
u- jt����Ԍ�x@�y_'��;��YM0OO.������Q1c���E�V�>�? Қ3{8�"�8����L�ݿ0�J� ����HF�D�}�A�"�L��,������bQx�NO5m��?��q��x��ho]�;������ ���`����i�f�GwK��O�uV����ڲ}^ъZ�>2��W��Hu�`j����?�������uU&u���u�cBB	v�	��s�^ɜ*��!�y��b����#�ü5��ޠ����W}49j�It>��$ޟ�4����	Go�\��t����~���P���0n�|�n�*����Qp�٭�Ƒ˺��=�1�&Y��{�	k-�X�����H�o�-�e���diHAD�9^�8;O��һ�W�3y��*Pc9��iN�&NN^��.�'쾉�Xp�r�yK�'�S�_�n�:L��P!��#�(%w4�)jf����҉����Lz�d%Έ�6KT����y��I��A�௓]��NF��?T�)���o��bwM�	eXc3D�v?kc��������	�xpQ�||�� k�4H��h���{���I��Pcr��C��tֶV��n�=�W.��8,H@O�;�z�#�F��'}��@�dM{֧O 8�ө}��GB��|��*5�iI�u�B+K�ЦW��T�֐��d��)�i@��u����ǽ{�%���XL��;V}���OuI4#|f�b���G�T�7<���`������+��#�N�x)�������1�B����".����Zy�6�/Ga8�؟�f���f
�-�E�0�o�<R�w��ɝ��u����C������S%BUmJ`ؼs�X/Ǹ�<�verw�9��-H�P�|Ҋ��M�/@�S�{|�(@~�I�m�QI�M���Hy2�¨n���ʠ���(����E����'�*$����c�"�G�tw����e6C�%v)�oޔqj=���>p3����hJ�B�T�qH�� �����w2QX0~B�ˋ���j(�LJ�&��xE�i1OE)�;XG�i��C�_�H���5���%7߅�|D&� �jʜ�s�V�s1.2��#�O��l��:Y��#)X�ۏ����^�l�7 ܵ�����	�ZKsL��("��+|�t���e7�=^������L��z>��<���&����+��Nzk.;�e�:�^=�^I�˩5� >��4(O��{5���7��{%r�<EP��U��3o3��~��+��h.+�r
"��e	5�|
��5*҉��O;�Y�,ߓ��z�o���|Vjd�����o_�пc�^��,O��75��"`n��gz[�N��Q.{�@Z�Ίԍ=,b2��2��9CD�m�s���ط�˙���Ͻ��{��뵡���O��"�j�?����|F���Z�]�Vj|G8}�C�?�y�~0�����urpȣ�<��=Gz�Ma�r��ɚ� �4.a��&�C�_e���e/󱐌�_��,*�ɷ��Fx�F�J6bP,`��c���Uu T�(�[)V ��e�^����&�9�Up���7
��&JJr�9���Mp;�=G����Uq�v��eR�e771��b����i��
[��W�߫�?��i�6<lh��"��߻���w��a����h�	M[a�� q`��L6�ɯ�T)�����$c��$�X��#�`rR	���n
���G��ϓ�{�j����������񝇊�o�k��~�tY�*�	t�h&/;;4;Oz	R�,J�Jk����*3]LM��[iC#��}�F���`�aќ�����l�-�;�r\�bY�mn���b�w�H�*�b��f���VE~�6�s��R3T����PA{q��䪤�.�6���ꋶ+��M*�A$�=� %��#T�r[1�>ة��A��������ڍW�%��b�Q5�ggζ��[GT��%���M���h��q	�]��;PZfX�b�J[G	aW�Ԗ�A���6K��u	T���^��K����HI��!9�Ւ	�2Ȱ8U�}��jzdԢ���*.��nu���:���b�Ǯ��s�H�sn���#A����1"��wG~�7[i�2��p�]\��q�����e��wQ�R"��<�.�Y7��i� &�Z=��cz�a�$�J�n��f4�jCb#�ʽ���J{<'?��ԙ�D��#��Cu@��
c���5�� 6L]}�
��ǹqQ���|Pp���O Z�d�z0�����Vv�dem�q�+�Z�v-)V'Q��\g!?}��L�Z�t���~ ֽ���y�H''÷�k>�,T
��B�Y�MIR�����x����gAzca �����h{ �k�mR�H�IL�>�>�03�NɃ@B$�Zr!u�|�oJ��ϲ�z���Z�O֪�ZQ���=������SW��EObi�0bin�DD���'�x�+~Xӻ���{�'	�M>��b��"�����r���o�.����� ����7�V-F��,l�1����}g�6i;/�!ˍ�B�7�#Q_Qђ9�Ŀ��bN�Q����P׽�^�vo5p^�� ����M�������@p�"�)�߮7�=UO��*/a,z#muRu�5ϝ>��?Sb���ls�<�W��g
�(!W>N�R������3�u$-l_�:�D�F�p|dļ�e�7 <��B`��C�7�և7�'�駝���c������N~�<n���T��)nv"*��q��`�p����1�� 
A�E�X�Fj�E/�;�X���>c�)�e�h�nfθ,�gH�-��@�UyVY��� �����z�njKݡ��� [����q�~M^^]�7��/�<�㒖��&����
X�A��
% �a�#"6Y�����|[����7r�gβ��V?��F���ǥ�5MG��/��7��%����'%���|�EE�����v�� ��x��S2�ps�O�&�n�����;Q+�ݪ����r�؂�z�\����)9�d�|�kd��[���o���M5�y��hZ(mU�{���"���Vod%����`t�E��'eH�J��v����G�h�E3y�$Z��i�N
b��n�.;��̟>���PU�k&�ل�	�+���c�}??�˗��?�t�1鍾"�mm�������;�P ������
ğ��j���(C�:����J	�0��$P�\��t����ԙXV�q��뫂l���t�̿�v�tm�<���u�ģ�/)�����l�C��d�s�؀Q�mhi	�,h[+"�}��ң='�[��-���u��#���K���dL����j|X����� o�
'�7ߑq�o���<���A��\�aaDS+Z��=n)W��������J�b���U]��fH������~Csj�_�Z�nɯ�̓�}�HFG��h�'�n��w�DZSg�̈́�I��3�s�D���D��Y�v_r-���ȍ_��@�F�xn|h2���f�)Ĕ�k���S�m�ҬFIR��2�Kj�	$�CL�Y,��M(Ɇ���q�Op>��QH$'%大�����������KH{�l�i�����dm���M�t����b�*�u`�o���(��N�L+�O��u�A9X�9�B�11�d�1ƞ�ᰬ�
9�� �B�0��қ����X�X9�������Ⴙ؏�ۻ��b#�&VVb'�8gS�Ft[�x̾a�H������Jg辱o3ԁZ�_��%^n���N 2��j0�}�G����Q��]�u�Ժ��X�?�?�>&iFAäG��[�B`*d�i�����DKγy	ʎ��.�2����(*�ԧ_��aa���%>��/٩�8}RL�HK$dBY�!Q�j�1�:o[G�X\o௬��k�{������_5[����xB�	���]�T�#uQ��7��
9Z����QRǲϒ!T�7��Q�&6�o@w���(�z_�����=�Y/k��U����h{&(�^�;qI)c��܀��_T�p*R���`�����3yu�BuW��CBy� �'�eO�>$$�1�:�]�C[��_^�t�~�6�O�*�rT�F����ńA���
���5̈��6�w���A�>��RD�(W'x����IxS�x�-J�HҾ��)C����)��닉�k{�T=&>7��`��N�)��O��9(�VW�>�>�O���7s�h��I�l-^D��=뉨�(�~:\_�z	2�����6`��oQ�>�����rH���tKȿċ+��&���ƍ>��=���[��S�W�@�7�et������wΊ�p���>a!�0 5Z~�޷�Y'�$��`J��K/�����}n�R��6.��q�<|гU&�d���� �f�Ρ�F	p&��j��e�*��t'�d��_[��嗻C��H��"̃3T�u;���i�M8�B,��:��ji@�qn��b-�bq4F�Gl�kD����&'5tR�й�?T����9P1���܎���	ed��V4(5�[8��U�s�t�&��Y5�������@3]���;��U�V��zw��@��!Q\Y���q�?��޹/(�
4�<Mn��:1��0�oϳ���Q؆�������M{�F	ѣ �����ɣ`[d��.�ڂ0�l	)��ި�s���ūu&������a���r�I$�q����'�h5~��&��¨.8>�Jc���a�'�oE2#j�����"#S�ܜ�4JW���y�a�j����2eU����1<.J�8q�]�~����YS������q3F��A(L'���:��Wb����kFt����=b~�#��C�%(VĻ���q��g�4^O!A��\(�}+�X� �c�m�-)�uY���l������t��g��9���'.S�b*����M2!��d�G=��x����)�[��� wj��=	T(sֆ��6�ͻ�2S��MS�~Kym�������5{|�hv�n����c��~el�kt���[���U2!JX����}�k\��B/�B;:�%fr����E����+E|��~}"��V89���yN�W�㢹q��p��i���Zf�O��J<㹤Iy�c ����t'/�7J�GQ������~�k�1���;�·�0�ww�JkIΉژ/��X�3��ߛi��F-͙!�>�����I�O�t�,"��i�2�?J&����y��.��_7
����Z��#*tǯ�n���d�+(.�>��W�ϱ�#��x����/x(5��e��N�L�؃Z�*��yTQF�^���+��d��c���t!?�؆!�����.��R��q3#c(�A�P}T���8�YÙ㭝}���u7�vw��X�OF֗D˯zRU]�J2�����	.�k�����7��d,܄��]B �7��q�4{<ݬ�X$>�9Ua�:�N�`N�K�Nx�_���&Į�f7nP.M��p���B����pJ��@���!M�� 	��9������d�h��`}p�xr�P�ռw����y��^�-D%q}����QRH�ӈ��z��C(�b�B/� �����p�r�=���g}f�M�{�9jp�R%'FW9h�@�DF>>��˽Pu������H���li��L�b3���*/�,=�{c'�ؽD-ë,"�cS]��^F�ֱ�|�+Ц��Ih2m�����y�����h���,�� �w^��(��r��B�fz�\�X��3�N�B^��dH�����!F��k��z�l�Ǆ��R�ﴌ��"��ja���U�_��}�Z0��͖0���Mc��˙^{o�j(��۵��А�GJ�6b��������*Q���E� &.��'u%���7���c؏�vv/�ɔ/�/�|�O��ws ��6갇x���՛�����d*�[��%�D�]u�]nnb�U���I���a���hz��D?���4�eܨ�YyɃ����OdˋriΪ ~��~�{��I�B4� �wE.�40�/����m���kܿ��S&Xw�F-��hKM�a<p��W"Ȧ^���"�}����1�ReT�B
�w��]h'>}������io�����"\�W���M��[�n�˅�l}��r�`�]��߹;�	,E��E�O<����\���Q�sC�ĺ"������_�l�fA�Un�qj��Uf��In�Q�� �U��WP0a��^�}<�p,s�V�	��QN�:��f1C�DV6̫W-����(+�,�������*��>s�W:ȉ���?\�I�� �j���NA�D��¼_���٨�-�TJ� 7w�L��jWey�Ue�D�g�d
~c�=M��8H�J`��o9����XF&Y�x�x'�he�㴾�;��"-��z����|R(}=JY�<O%�0�ׅ��m�V�� Z2Oy��^�ӸnZ����vQ�j���ǳ��=ߍ��p��?��r�t���ӝH��/::�7��6U�) �5�t0�fD4�p�{�N��h�P����Um���vV�0���}������])���5T��<.��XRL�wZ�l��^�ܻl�\<uu��hX�J@��aV&���9�ql���O�	\�:�vMM͚��@���䆸�t4xW��~5�{^��\Y�����X��l�LH�R�ꂡK�07_��$2��N�|��J��N�l0�t�Ib#��p�۵�o7��8Ml�y͟�b��z��VT�:�k!:q%��خr^��4q/�17�f����v�WB��#)&�ݡWj�/P|Ȫ�E�E�]��0���I������ʢ�0�_�h
<A����]�`�S��K!�V8uB?@^�����\Mڶy�m~^IHi��J
�����r�(�|fHt�5HR�,�	��Y'ʖ�$��ՓhS��9�ݹ�6��C�ψ��М�5���.��4#Z�L1��e�`�l5�r���C'��yB;�>׫�م*�s5~sH8N�b�W{�O(�ƿ��jD0����ݚ�c��׊e���t�k�������8��Q/�z��vRkk]�����7ߍ�/�&����Q�HY�x��J�g�Y
h���b��Y��s�5q_��7g� r��������(t5�|�@\/ �Y�o'�7e�s4h�'y�Fߛ��as]RXK����>o��B��k�"���2T�� ����/��t����P؎d��{IHx)�H��mYm�p��c���[ګ�sj���dnwP0�M���M
��<��¨�c���6�H���dm�Od�����kA.c�T�7o��x�p��E6N�Ş�)V�'x�E�p�����-����1l�a�t�.kS�ܦ���^�~�!��� d��L@�ߏm�c�R��^[�#����|�;֕�G˚Y�Ϗ��	�vP�GG��F�����O`���Ӕ�]�͓��NMO7����i-.�s��cǒ��^�@��{
!N����-)as��Ň� \ ���M�u����O0CF�)i�>_�Ul^ao�����Kl�*l�艤/�۶W����&�LT��O���n��Sx��YYw�{������7{�g�:\]��Qk�;L��=K!4�����5�[[����1�z�_��3K}S����Žá;��	�g��8Ǆ��_��/2�����ꨨ���CRJJ�")�-�(�݈t���3��"-!)� 9�    �� 9� C|g���~k}���z]�9{��y��y�~�9>�B�PE�/��~����B��z6=��[������YcAHZFPE+���m�3_���}/N��ɮ��G%FUY����͎Q̡��̈����GS
�7s�&Q�p�Є{�ڢ;p:�d�J����� ��U������>�V��ރ�eȢ����_fF`⧵����}�o�7&W�RF�s���8UJ"�e��yw�׳b�����i@�WL}�P�0���;��(2�8q"I�hR{��y��-t��P<m����BWUi���W$�����s_��-�}�<��jb�����Ź���\�h�OO
D�t���S�T���^S�W�eˁ��7jxnV�z�r������ؿ�m�k
%�=`�u@2���F~����aBʞ��7I�Nc���pP^�|F	����C�~���R[SWr|��3d�rN�.�J05�67w���R ��X����n���`����q���F���@�C��<�1Uk��?�|�ϓX1 ���M�7�=��k�\�o��>��r������M ��wk�0�����%��f=�pA_H#wO�p#����ވ�+k�(X�,O%%�p,��R_�c���׮vq�Q�Sc���*���x�x^��.�P%��41W�SE3���ƪ� �|V�|6�=��E&j$.����j�`a���z~�
��t��0l��))���x�Dk�T����k� M�ب�|{��<�	�%��J���&�~�H~u�{T�6�@F���u�c;Rgɮ�:i���Ղ���Ћ߼�pY��9o�o� ��Iɚn�UEg��Ǌ`�������f�����!I��T ��oë��bT0��b�Z�ݪ�}ӎ����s9�#klbB	w���d��y�'Qm�&)���/D훹�/���;*���k��w�0�����Վ\�.�k��.ڴ������ݥ*RB�<�@y�|`�����pa"�v��r��Y��������-X��I��z��m\�� �zgY9gJո#{�eE����*zi�G���:b����j�'!,i�p�K�8st)���.����H�-��E�� ?�9���r��x[ٺ���g>�l�k��t�u��O��l>�%|�W�j���lN�6�E�������i�i������K���c  ɞ��"�.�"{�Ȗ;�[���
����K8�/�����0ֶ��4j4<�M{;��)��# �Mb���~4�����`fe�nQZ�B�;�����:8�}^Q�[+b\.E��qN��k
��B����冣�\����-P��衽��r����B�:z.L�N����t���H�d���������#UN:>u����ą�=e]H����5�?7�p��Wa��`�r���R�Q�
;�x�L�SO��0BO��W�'�XXb��q~��#�~����`~Fێ�:m�.��T�*C�t
?��t6.�S��	���=��+#�q��F��`^�w��;�cj�s�;�`ȷj���֔��������oQ���o.椒��ZS���tL�9%u���_
�������<$�t&��)з ��yƯ�E��#7�j�0N#�sr�p��c�+����=*�Q��>��Rn�G���)�N��g�HY6S�Q��66lB��D�m�Kd&6)��'���YcaG\�~��A8�����9pu�5;��F.��j����w1�=L"��C���&cB��@��ZQ������-��$
"��y4��]�T`Y�����Zh��ځ�g�ô�LBɢ؄D��VY��r����y��w".�5x�1FUo�T|8�tLLrr|�zst`��1��SI��i���;��$^\^��� )R�C�%z��1U�&T&*�=�BW���6���k|T�l�Fn��
N�L�zg+��'�*ѝ���$<eB|�2�O����bK!�:Ĩ�WnOm=�����nɊ��5j�B~������v}ĈOt�vg�p�颫��iCa������0�3Ά���g	�џ��5~ĳ���7����t�"ID/M6��a$N�p�.��|��
Bl$���\1t$�L�!����	I�� b�{Z�>��ό�eX-�U��H���L����&8������	�<y����˅�S⻨����oڧ�t�� ����vt��#m}R���oB"�I�����{����JJc�ՁgV����|�O�%9m�q���8�k]f��Y"�
j>˰�ֲ�W$TV�*��^��)����I��b#��ސ�~�����Ol+���O���n~�L�74U���$�����ʫ���O�����|�*�[D��i�z��q�o�3���,c��#"O����/������vʖ+@�
bIket�������qZǙ���J��j8�j�-gF�Vl^(���ߗKJ)�t���]X؊�WJ, -��WѾwo�+��3s[lJL�z<>1n�1������gCw�tf�̆W�@����~I��t�_�nn��.辵� ���q�cĞ
�h�TQN��~�^4��x�}��S{�q��U����Q�U|ٱ��Wh��g}F�Zh�-����ܒv�Q��0�m|?�����g�Ʉ=9�͢��Nl���eˑ@�}����J;�~l�6qˋvdf� &4��J�+zä�S��ۻë��|���l��������u�$��%�����2����[����s��JDH�p�����Wǁ�ǧ�g2�)���% ����w�`*�5��j�*-����k����ӊ�?�lH��lU���ϐ����O�T�%����n}Ya�"a�#+�C�T�嫇�-`�،y��/�	g��X�1 "�,ʼPP����J����u�1�zd&u��]����95���Q�,�w��7/f��~'ݎ���b�a^���͒�.�>l^�n��Ȭ�fnO�E�z�A��2/<�	p���{EA蹌)Ɉ�c ɨ����O����k����/�*!�+XRĴ�'�NOFn�E=ÞbtC����ǘ���J�ts�5K�*�����CeR����XJEt(mgm��u}q�����Ug��
�;z�8N�9���{{Ka���>�ۺ��7|����d0D��HI�o�PM�N�M���]�L�o����Ѽ�nt�@{\I�'�Y�/�a��w�_E��Ȟ����_�B�5]�b���xf�h�;���Y��a���5ܴ�g��v5�'8���w�#��E-Y�	��WU�{��h�M���UQa��#5�F[����A�n�N���	F '����:����&�y��.\��0Hlr>�il^֮o�Wݒj��Lm�pf��n��A�U��d��שDad�2����Z�Jg��{ڣ���As0�;�zy�_���:�6���ɦ�5r|�B��#�<��$�m��&����K^�rYЌ�#�!y���f�Nɝ�tT�A\s�uּ�z	K����ȸ��ۉX�>�ӏLJ?�aS�P�j�&��^s�/��*�N��D6�w�v�]$��YŮ'G�����J�T^��)l�X�=2ʢ�u����*���VDm�	�{��gi���#+I�B���UE1���l�r�A���#w:['�ϼ�K�޾&��d������ϳ'������$��.{���/�}�9�C�S{�ZB�;g"�\�y��*����r1r�lC�@6��y�gX�����f�\)�q��ʹO�]%F�}|jW��1��ڒD�дZjY�`j���5����S�T}����ԀAU8�����?����΁3�=���w��W�j��sd)�7]��qT��b��HLJ�EE��}��I|�pÑ]'�b�_���.����PH�_�u{j׫"k}<��k8\})�'��U<p��������r�����(*��N�#�/�����th�*4n`���y	&,6��bVEa���$�u���w��N����ﯺT�2����w` a1"����������_ճ�,�=�t�1ޡr�=8��H�����t��Pj�N`�4�$��ǧү2�1�k���uS?cr�sw�ϫ�?�x��w��
"����~������z�Ycj��2/��)&2�'�
�'�L�Ʀ�����R�y��Z���3~��ձ��؈0�E[���8�֟���
����M��L�ݰ"s.�Ha�?̢�R/uNW�y�� ����Ͽd���t�n��6!�oRa�vR����\�Q�����9�n%�]w�Q�����M�Q�1m�
�1�-��5���ȿ�b�A���l_�F�ܵ���Q:u��n��o�Uc2�o�@Z�J�NB�����A�*��8���{8<�>��&�В�M��c��.?�B,g|߄�8,eN�}�X��X�?j������Ak~�o��a��"�X�{ ���`�������з���K_a�B��Rj�����f�yO$��; 
)VJy�C1�n��u���Rs� � ��ox���sb�u��E�b���ZC�O��N�{���22�)��,����(�~f��{Bʨ�M]6/Ɗ/�H쫐1��=�'K,��=���tv�q^���r�\, (�gIs�Ѩ�zF�eE���(B�ʖoV��P��HP��\w���-�r�6!�;8%���\Yg�g5:;���*��QD�$Dd ��@�,��l��[!����EIgf��ԝږMޝa,�0�/�в`V⊪ǽ��4�Yسb�z�+O�F��q���J�c�S.W�6���ΟL(�v��{ojwS�&m���F}{a���O�Ur$Ȟ�����E���1������%yr��1�����N�bN8�W^L$o�ǘT�����	�G�c�^Y��!!H3�Ca� �qz�|�W��o�+�;�U�:���w� l����͠{�����
 q�N{�q:����t�k��cf
"D依Ea��VU��z�	\ȑ�h1��1�ۻ�pnCja�_1�囱gO�G�L�<T���0q2�+�/9�V���$�$3�χ[]�7/y_�:F�FF�c�}d!/���z��r3}��vGg��z�ZA;r�Ǻ����[W�K5+^��zPT;鸬k��0������j��Y��l�c||�ar�:a�r����� VW���zaj��U2�̱
�=��|Ӭȼ�hb"�@�^�Fm�0��"��!��QR�bE�Mof�� ��l�5orB�W���6����I;�G�����zДx��
�{p�M���Xr��
�"u1C�]|Z��|9A�2�v���`�)1�-P.���	g�%K����g:X�ь�>,TU-˔������M�4[̭*�*,@2����ah�U�qؕc���ی�7&z�KiK��M<��8ڞE�t�=5H�E�|��d�0��y�-�W��s��{�6!�|��ˣ��� �p$����1 f�✦ �@J���J�����;*w�t�0T�=�wB�_�wڤ�I��7�R�z|>���� ǹ/���|�}�E�'t&5���l׏�������^^�x͇u�+l��U�y811��}�r
=��1���w�t-0TG<�7�9Ѓ���ic�`���>���S��`ⱖ$���u�Ԫ�0�xo��M��M*����^p�KH��;���{�L?�*���&q���h_)�V@�bǏ�2e�۸lc��K�Լk�[>[�>;m����9i0�r<j�K{U�6ѻ���bγ5�5�G�l5���ܤ��$� ��vh]��d��/��둪�� ��RXׇ읈��.��s�7�[��?��
M�ȍ���g��Aw�u�#�4�~g��Tk����>E�Ct�g�8G;�����c��x);�ɘ�������x��xV2Q�9�$u>(:��
��U� Y�NT�t~�r���F����@����H�@�^�_:���n9�;����L������ڈ�_��4�!o���KQ��|��しoUf!o�S����ӺeG�n����ӯH���t�����R;��QD�}��|��ba����/��#amȧ~�6�f���ӓq1ku��M��/�<MJ���:�.�Z��\s���͉��e�bַ���v�����H�g��n��ϲ��υk3J��#��`?������pw��.{XeTe1�zz�R��̢�@P�Jg��z�իN�\�b2Z��,�8�1_l�^�ϛ���wRBe�d�%��ѷRR�L���Ժ~�čǘ��x��kG��Q
�����+� ���8ʐ?/�M=)g���,<��@�Y��B��������r���ݶ�B&�Ю��WY��5ϳ�k�@-Կ�� r�N��bd�UN�Օ�c9e��>�U�S�M�G*�I�Ŏ����P/��k�䰟~8'$�:1��wRΫ���\\|���#�NkLo��������?;Sܬ�I)\ّ��Y����n��%����}�庡`
Z����S/��Qi��F_�z!�-�<�A˴wI�����s�S������l�6j�s����>��p&&
J3�W:M�$u�2�k-�cn�bO` �,���Sz�3�;�W-_�\�'6�i� ���x�s�F#�1�e3��:���y�s\1&M�`�Z�w|�n���m|{��ԗ�����P1O��N3��3�GR�Ľ���@�����1����ˏ���� <��AI�\m���b�}�K.�b�T�S��g���(;b�~~��>�;�����F��߶�����ep�MH����<j�l+5EI��{w�i�A�e���Qz���,�|(2_�0q��ycڌ'E[���+�U������{~��V_�u~L��(�]�+�����w�d����%���q'm��`�+^!q\���Գ�+��%*� ��Ə��/�N�Ο��i�=@gG9Gu� ��p]�5(�Z��Uߟ��©��é9�M��&i��g��3Ry/��w�f�v���[u�������A
����>	�]��+��g�|t#G�Tk�2�p��NQ5�_{��r8�H���=eװ��NՁ�23��q
�J���K�/�\=T[�!���T���tA��S6�bK$gr������J�y�b��F��k]�gj�
�o�d�#��HCcq�>��U��Ԑ�M��	
�������x��-m�|���^���kz�A�k�t��d���b
Bk��*������g���2~L%L��\����j����$�����H��!A�T�m�ϡ\[�z$L��J���\Tz�:Rc�����LƳ�+�lK�J ���3z�R(�>�,i�+\�SF��o�yD�\���=IZ�M)A�"V4�`~d�e=�Q�ŗ).�%������T_��Z�~�Z��d��"2�J��N�L�ю(��k����S� rașTy��R��z�l����Y*2AJd���tZ�(<[䓰G�i%�����N�N3�-p������]�@fD��l�ʣO|��v���� ܇����v�d��6����� �k��)���"��ba	�3�gr�Qҥ���1+���7�'�1z"YT$˾^
�ޗ�C��ֈ�77�%n;'���LHX�0�5����փ�#\��?2F��Ea�`�E<EE��8'���g�t���������|j�UCra�6�kNV���.S;/�#��'�������:���;�L����s�^h�b��ՕX���G����eϳ++�]Q�A��4@��	�:�ʟ)o���|H"�>m��A�I���,�^˖�[/���j8
�T"���/�|�$��͹��2ڏ�Y��Z?�;e��Qg��4�nT0�_%���w� Ỹ��u�Nc�%�^�r&Ϲ���i�|+�n^�G�)�&��b6�gԌ���Կ�7������9X~Ƌ�1�3ry�Mm��m��K��8O.�#�;n�4�tȇ]�:3.Nmߞ+x���� x�<��v&<�:����v�z�߁ؖk	��9�^]7�l�J\O;m��3�t7�;���vw�4�ţw�g[��7p�+���^�
<Co7ST�lix���$0Ya�(�F��X�D,<�S_��Uf�vA��i�B3�Po��H�/Z�����ŕ��-w��	,`��ԋ�J>.yfO3O�Y;y�zI��[0}گ�GU���^�80i*��[>*�/���+\� ����1P�l���ӥ������i��p���"ے6�П.����L�5]�t�� �6�<$n�)m�/c��)���G_���X�ߏ�w�:�=�m�d�'�.���������着D"��)h�<"�%���N��hh�Kq\.�ё��o�(�Z����䋞��mww�I�p��xֿw$`b'ӛ�6�o����4��t�Cb_5�j�F���N8A%=�h_p���5��-[V!��-Al3�ٍ+)��߆�gk�Qawvs�Bg~��'m��Mt������}�>�1�[0Zb@:00޸��p��d��ϲe� ������k?a9S��/��e&�����.>�)"�B�h{U�`e���k ��V��kk!��-�� M�Љ�cr �>%�z���o��j�����u��,��x��ͥ
�4J���n}v�v6/�ʎOw��,�u&� ��T�rd�;�	1�-������>��o$(��y�Vڨ@ޓϲ?����F��w\	r�{ LgMv0^��o5@ެ�\�����!*R��9�g�	��?LM	_3#�ƑKǧ#b�mz��y��ʀb�o�p�	=*�@����5/�c���ۓͥlS�	3�K.�7XS�ү�9���tTAhu,��lNԟR������n�;=Z���ÿ����R?��۫D�@�?bm� 966bB���aP���)E��_�!��f?[�X��{�S��e�u=7kB\��*�H�_%6�M����0���eS*�C@4�J�R����Q��B�1�9a��x ��i�
�ߡ�} MQ65E ���h��/��a��;����{�^"����΋�/㍅s��e9$	A�&�AM�UU����-|*<ch/��T~��K-����BoPT;D3'��O/vbq!��F�����M�BN/��Oo�O5��BG39v^Z<���������{<0��Lb �S���D�2��4NP�R��F�!$�j6%���R����<D�a����)5�Haӧ���?pvsT�M1�ФF=1U��B�5����ݣ����3(��HU��p
S�l�(�;o㎫�|�-�N��(��.����smT�NN����YK$[H�o>�m$��4A�C@+$��r��ﷀ80��44t$�wS&�����M7���Sl͔�k@��'�[�*O��0����6�G$D}�B���Ћ�^�����Ɲp�D�����4��$2z�W&��ZK����iX�G2<����%�!��m��@f�4����Ab�q?��6^��ז6 W��Hm�d�B�}�W{,�U�  W
�)�ץ��F���	�)H����C���DN�)���g~�
�n�r������K�zğ{V(�E�J+��[S$�;>�2ܤV�!��|�n�ǯu�20`��йR%�7O�J�<��vT������iEʷ[����gk�{
��<�{~�Ϯ�;�n���_]}��ߝ`L�W!ߧ����x� �L��yT��x�����w��n`�d]�U�r.���)k�tv��n��c�2ڏV� ��?�"5�6��:hŵ���q!��ԛQpp��
��[c�V9��G��cO���ߏ�ʎ0��[�ޫ�c}R�ȫ��Y_� F ���Ϫ���NA^�Թ��`�BtXA^�B�h����B��%����y�J�=��)쒱�r��"�[�9��1xt�r�wJ<�й��h�:���iW�p�9���YU�A����t��ªc�����?����p�Y�w���S�e��i��t���3�>�q��f�-8/q�����S�zl�.��"7�jEF��K��#��+��}�>ݜ9��t�6R�J�ݷ{�����Rqg�'w���@K�{.�@h��sr^�`aBf�&N~+(�[����P�����c�\��{12�H
��@�j7�������i_RO�)�̆y�=
��)��Y`��[{sO�(�O�X�%#F�6��آڟ.C@B��
��cMZ
��#3s|P���	8M���VXOʐ��^�;\�Ь�$�8�ͷ�"uʮh���z�>5�/��ه\~�e~_�q_����z���?��<PDۈ-��EvR'���\8}@���,n�_X���ߪ7`���m��v��/���n�ߴ�d)u�_�EU_D�����Y=��ˑ�X�c�u�}s��H�t<72�p��V�X�u���p9����9hu���� �M&�p|iȝ)o���`�Zտ�DR��`��Z8́v	�mkj+=r�q0�Y�<P��h��Ňp�m	��d,Q'�[SΈ�s�"��}I�����%�d����D��S�>�.F!ї�����'�\���@��p�̥�&A�GV�kkA�Ʒ�o����&$�I�H5^oo�ET��K4��q�7�nKmѓ-�n�p��8X9�k6��yi��h7w��?�i�ЙKy���Kr	��[Q�-��m�_�B��Fz}#������� ۫���A������ܕ��>�_RJhb�iȏ������VP{6J�+0/�__�O��f��Y������&���"��cw��I�>o��HШ�ۋ���Eɕ��H�j)��6*哤&ѵ�`/��1���):�y�yW�p9�����e6�z��GM��y��S�ͨ���,J�(7���[���ۿ�-�iͺ��V�BrU�G�VΝz ʴ�w+y�CZ}ՏQ�W��+��O�ߌ����CPQ1���D�3�aX�ۤΌ�Y���زd;ܠ$�(%
�92&n�e �OHv�tNT����r��h͐�ԓ��x�`_��P�Ḕ�1����*����` A�)>[z�#�g�#c	��^-+Z jd�,�� j5���L�H=A��]�'k@l[���a� roW�����н���i4"��Ƽ�g0.�w�&r��) �E#%��69o2��u�画0��-H4!}Ɯ[��L`��/���[p�ap�,�L�lX��b8#c����ZV�I��x��Q��Ol��Hl-�%$�_`�}���ܬ�X�y������硔ܾ��~W���c����'5��ӭXV��}���$�^��~��>�-$�=I�2.�Oy�^$ KE:OF��'ٵc �5��2�@܉ޏ�Ы�fm;�����T�mH$u�S�y�ү�S�|�Q!|-^�`Cb@.�O�~օQ�΅��\n�ն�!��� ~ H�����G_Z�/�,�^��M�3���#�g:S�WЋ�#�#gp���1)2��������`�Y�L!�����;��ͮv�ՙѮ��4���!�cD��Cy�h��/�E�a�L��b 9H�c!��=���n���e�юq��l)��5���������􏩃Ǻ���b3�@_���?i�������Z�xR�����R�w�>�c"���(�U.��푒&��.ZA�1qD��;
h-8�V�$�6!;�f��O[-�<-:�ͫ��\�g�ƒ�a�<]7	&X:����^<��{����{tBfq�eM0Ú땄f&*�TW�u�?� ��R��8�F���mL[�67t=�n��cN�����D����� �-yQ"8w+�y ��H7��^GN/�@&��emS�	r���J��mU��x�o������ ��o�s�W���	���qaP�c�� -Fn2��ꍚR;����ށޔ<j�W�4OL�HLZ
�������b�j�b�ni~ΰ�3���2�\l��l���[�J���۪C����H];�;��  ���AWװvWڗ����%�]|�3�����^�][T�v��7���_j�Q'�g.�3p����9��v ��;5��'����oIo���ؔ@�14��ǿ;B��i-O��ׯ����X���3��z�Й����]��p������$��3�^�{"|����j�[i�3?g��;���o*��"�م����U%%R������6�nc`x����IÌH�ו﷈wHpo%�O�@��Ҕ�� D�;V�.d�C�%��� ���dŗ���Q���f��7�<�6���ʣ��-�5��]P�jgD�K(�7�r*ͥ���z�}��zc�׌�����R����p�x�!AD�=���Y��r�Z�ٶ� ��г���"�32ğ���Y�j����)#� ����'��ک�#�G�x���~�!��]Q>�7L���̣J�`����:*�'��OM���-��çV�.8�#Y�Kϟ��[��_'m0�V&`���?j�,����ro�f3t�]��?dz�o�aO���Y�V±r��h�	�;�1p9�֜��%��&�()�e��?����.��j�+�"D����X���P�8|A�0%娆 ��#c5��%W�v�%���&gZ�+�H�q�� �e�[5��%I!������P>2gĜ-d6��1��C�;K�JsK4:��Oho_x�m����q��afv�#X�O�ٟ��m���U��)�I����Q�/��`o^e��y����5�\�������; �������P�E���Ku�ׂ�nхsa�t����0�ސJ>5f���.n�N�֐$ :��셈�*\��x���L8�Z`Ϛׇ��9��2ľ[{��<܇��2��07�:%��T��Y�G�fR��.��ES\���B�Qh툉��EI�痧���»���m!r0���R��iu�ϛ��q�@7�pd�q�ФQ@`&�j
!|��*j������Ǯ�����u�V����r̲<<��Hۚ8�O`��{t�#�85��/��ǉ�8��A����=_���1/׳pj�:O�� |s��o�d�.�^���77��&+Z���SJ�ƴ���J���N�W�R��z����''�O�X��P'A���n�۩�Z7��<^a��I���lU�����k:���*��Ȟ����P��=����Nj��GZ�A��cՀH8�=ݍ�QBb�Ao��L��cp�X��EY�.��=Ø�g>��O8���L��l�`�	���${BW�����Kw}D�kZ��<+]�Nυ���;]!["�Ϡ��B@��:�|聘xE���+)NA�r(�s�=58��1-[!�Ng���1 H�'��|)�M�����?�b����YSN�����1�vEx�sP.��sPZ��x������ssm�l����`������xr�o-8�<l�ɦ�}{W��LX�X�l,(9突:�o�6����#��kF�R�����q��"�r��2��	�h)!5�!�" Of�&y�� ���\���V����kd^z��h������A�OK&�B�x�k�A�%)���C�N:[���A�1}H)MG���z��X#K(<o�c�����ж������0qՉB�?�[^����@rYT��Gc)u�-3_η[%�F$=�����s7߹��զ�]��n���q�:�u��E&X��|ď�k��*��B��>8#[ջ�1&$$�;6�"�.a	���
2���kO��ft"��fe�~4MS�S{9j��;�����bn�J�M`9����r�}��#�+i.]�����>��KJ%4�ZJ�?C�1���QT��@��>�l3�~��!XO�o`
r���������Q������|d�2�x�����(�6��V��n?���
y9�F��"g����΁-x�q'�B�}��烳��C��HA�������F�z VAΥ[�4�#)�����at��@YT���������c����f�G��vD�b�����xI�`�[�4�i|��x�{�;����U������kC�Ho��FNj�������6@*�"y\��U�;��4��Z����i�g�N�oJ4	H5�"m�,MG/��^����^����v8��~4�s�tL\^ϔE@O=./p ��67����=���p!Gߞ�ҹ�z�N��Np�i�R�5��)�5���#�fC����uǅ4��ʈ;y��]��s�0\�n�܅Dbp�u
a����Op�9c�P�����@����p���⁹�K�Ƭ'NꍷF�����V��,i���X��`\��rj�;3�W]vU��*? ^=�����T�����F"�ޒv�z_����DrX?�>V�����5o���~�&p�����Aߺ�'R��p�"gL��gB�.o(��_i�<bM���F���B����]�]Ӯ���o�X1᫸�LD�V�+������R�__�wq�U]�I�2BB)+�{R�<�Μ��]�x]�H�nBm]�����{�ɮr�h����X��H��ľgƀ��<��,Ϛ���R!��+X��Y�d�9|eG���s�K>!ê��8
N�k��-�� Ζ�󭬞�����Q��1g	.�R�l�*��Z�U»��� ��a�&Xv_Y
���|��&Vĩ0O�Bg��Gf����GD�像�Boj8��8単4�J�͋��L��)����3�=��,Kd���=����_�m�Ʉ������H�_�"��:�p�y������c��{Gk:tՊ_ޞ�"�#��)����M�{V~HZ��׋X�Az,Hl��1c�߱���If�G�3C�t.Ժ�U$�7���͖(��ԈI���8��$��8f��ԗ��_�(��|~����e�OG�Eo$�e�A�̼�hs�&0f��pF\\k gq��t+	��J������0+wA��@�]��h�s/F��0a�8�2�R�-j�e�X����x�ѽ�	TnՐ��z��D���w.��rR��L-����@�ĳA�͆����o��]E�Y)��1��".�t%���c��4�b��0����4��8��"�rpvt$��'%��`������_�:��#�J��V.�nY�������N�q�?��L�7�P-I�`B`�N�:~l�,�F伡.����#�͠ �Ws�|``5幰�])��f��Ø���t�&u`�4S ���U�����}6�7��Ō����*�G���Ƿ�rᓭ)~V�'3 �"�F�0����Չ���@
70���~ȞJZ���j�${f/2V�xﲨX��j~d~��_�5ԭ��΃�@�;�^�#��|��bs����/�����B_r����;.h��v�����7�\��T�$Y��I�Ĳk�[����D;����2�N��ͳ� �u�՘gAg?R��t�̲?�/H����_}-�U郎�\���S���*��.�w�K�հ��쨣�ѷY� ���Nɱ��4}�b���~i-/�d�^�Qͣ�(uv��39E� �����5�6`�y�\���P���+�i����??	'�IP�M�����涚�eּ��,P��ޫ���?c����;�T������z�v� ����D�pך���x˙sy����mb��O�<��i��>j�	&�y�^�N�بgk���$�t��7r��J���\��\�յ��KK�
M�{33MPT�<>^���@�ۯp� ����%�vf[�)偝Ebb��o�ž�Vb��̏��W�\}�B&�'+�Bx�a���Ow�Ծ��o,�������M����G4���
ڝ�������_0G�����"��<�Q�w}g�Py��?�ž�h�sM�z� )\��<!l��B�װl>�z��PJ;\*r�ߋRk:?�����3��	Zm
{�7�1?����̱ٙ�ة�LtM��[?I�/h�W�jI���@�u�;�5Ew�z
�^�� ��S.}%M�6�)9�w��}��$����o΍F���LW�� �L�zń^z���P�q�⺵ԕ�+H�Ry���@�[>��Gv�L[�(�g��;q����?R�G
X�-zE!^>�K�������{�k�q����%e�1�4�Q��h�k�;��A�:�pb��l�8�8dH+UM�O{���8(��sb�G;b�N]�o�l���>�?]�[���]�I�(��Em ��i��G�\���uc#����U�F}�����b�i�Q�>	H҈ɅA����
*�O.<|�f����������8WZ����2s�^��ptzt��xؒ��/'cY��z�$���x��\�����嶐�G=u�A��)�����A���oȵ��5����]�7�
�.a!��X�N�I�{��t?�K�;;x�hg7}��2ᐺǸ��ׯ&�]�oG�Q7�v]�ŴG�%�U�i�{Vjp������xD��u�ErvR�Y�� `?AHid�,�� R�~�I]5� wEu)����^�u^I��V���RHFM��r�R_j_�-jyOW��U�k��W��+��5�=���X�l@����ۏ�1�J�C�o������a��l��d���l`�B�{-V+;�
��L��5��C�3愴����Q�W" L5EŽݘ��U��w�/�%�4_Y1��s%7ކ�R���0�I��^V�L�Cu{*�v� �g�+��w����3� !�� �c�n�r��
e�ـ]m��m�Kx�ir��Ŀ����%��`�#�@,�G�!��tEvYd�p'_2yh8�q�q�����HA�P�����tF]@zgΦ���g��&,��ס������2�i�t�L������mt���x��$n"CsO�e��!x��CWdU���C�Ψu+���u��%.��8�7m�i�4ҿ�g��<�)����l�o$�����K��a ]�����P��t�X��2��q���*S+��]���m7����S�&�'��8^��Q/��x�1<,S<�>T�5�^>�&J�k|̻�ru2����m<�2{�ǃ����mR�-���Gq�{ܼ�������z�޽�%4=[�[98�h��W4�����'����f���U�.O�%�6�4�56tL�}�n%� �̶����m�%2��筰3�uX=�$����k��iJ��H��ۏ����V�z������:�3)y���$^9��g�x���Q �3�;�3�#F��΍�f�4^�;5G��;k9%&�> y�#�h\����B��W�}N=tx��
ĩ�Dj���
qa��&���D�����aM�]�p\��Ea]�""J�^�G���ґ�Kh��(u�5�D@@@zOP�K�:��BK��L�}�x��}?���t23gN��}��Mfr��2�Tl��zΉ}^�S�j6�u2alr�2�X˕#��������L���'�t�@�n�ʀ���iq���@>Z9N@�3���6��h?'�Ӯ&a��H�O	����a|gO��\E����ʇ�q8X�9���*�R������ӐC�1ev�)����4�X�o�9�K	���!
+�WoO�l~"|:?p�s��Y�ȫJ�{�4��yz2+��^WA�
eQg���K�wE�V�Q7����sH�._-'��/ �^\�5�󹾯r��v�yN�>{��M����Ҍ1?Y��X��"2}[�~�ҭ=��t��f�D`a���՜��l.��-s\QY$�KJF�٢�ܲ7j�Y�����8���*��]��zz�.�yM����=����tqV�����v-���x�{6Z��ʗ�̝V}�A:�OfV��>yf�c��5Bz]jm:��ܹ��|k�Z㽫�n�� $>}"u����m�����pFf&�;6p�����Ȍ�{%�2�&8��!���a>������R�c�Jv6Jv�dg��Hֵ��d����3[U�`(�gȔ�����������fz�� Y�E���N<CS����=0���s��~���q��ʵ��Y?\i�u�w�*�8`溯8��`�K�M��ޭqT��᪡/�u&]l_A�X���e|Y_=i2Ns��i�������Hc<�n�t]��K�Z�3��9�;6��ǳ�'>��:χ�,+��ȶ0�~"2�8��:.��R-�2�Z�#��|��ҋ���+�o��6��l�>/�Ђ�w��,��}�A�@�!�xb���c0+$��:�8�Y���~����1�=-�V	���w����%u Yx{M<�2�j%W}�{:�1���d9��$ĕ�X#��²��:+��I���B�</8��Ռ����ȸ���y� r�O1��d��؜�L���fzg�~W��,݁>&�~z���#^�5G֐�[���#6{7]^N� ���w�Vp3�X��Tr�Oʫ����z�Z#95kē
0�镃�	?�78P�==��W��3us7�I�ە�Z��?qM�"_��H�O�e{�0f�t�bf�`f�����pn�����/E��?�e��z�I�f���wŗ�@:��N�r�H#�2�TJG�|X��R�O��!��@l�h8`�BL��e�vC��Yi�/޺y*n��)t-��₨G@�1�1r�������~�ͣ�1��n[��Vz��T&7 M�o�2fr2f��4O?��҃<��*k�j�D�Ʒ�_)�?�E����B�?m����z�x�TNn��i�N+p��%��m��X�>��B��`oq��T��l��F�nL�6��N�ʗ{�Én���_WۡBPg�����6i堾e�s��#e�Yj������E|�*m���4G��ϫ-��;�$�;p¯[����ٗT%���c�%��P"�"cNwbp��K�����(���E=��]8O\�������������嶟��K��b���.�7�����n�j޽k��Ok����������S��oz��jߛ6x��X@?���t��E9b�3��Ҏ�������S����� 4�}�]�7��B��A��6+�&�О�[��] 4��；��c�T���ESx�
��
{����Ș�Y�l�3�Uos���w:�^@";S�k�q�쾮@�X^dK�OAt�����]7�(Μ:����C
B��ʧM���)�a�����Y� ��
b�5�j�8�	�	�SW��C���� ��Z��^�b���•�L˽��S�N��'/ĝ8s{j�	�25z�O� ��3VR�������G���@J��:ޯ/g0Z�'�4��*܍)�`�EY�`��?3��-'�k7N�66�)�z�uQqϯ��"���2���ϳ.�}�d��e**EV��	� ��t* C�W�$a7R_<�#!Z��w��l\]I�g�	a����o�@J�X�vXLt��R~����n-k�_?w��K5X�_����c��>dx!�R/�qt���%��ޢ9crc��r��������ڧ�/Zj��|��"U�g����"�m�%Wֶ?�nw���x�v_��.@T��J�?�ܟC��:����3�ţ�|�Ej�F��#d[�孏�|N1���,�v���gw�l��!�<ǀA�[�=�9m3��Q;ϙ�G�f���u���A�|m���;=wý����3`�5��`#�qO6���_r7��}()��cOm'��NO|���?���U�滥fvZ��%�1���� �Al@�  J�����t�5o��V� �˕6p:���Ѽ���!��O!V]�jN9m�� 4m5S�FE���J�/�*���̖����n?���Q.��kk̛�~ԝ�H�Z�����b_N2�^엻�"#)Ȟ��p�˷��F��>�x��	�ష����u���R�(6O?��7��+�����L��Ypv��*/gcO�O�kU'�UY�����U���2ڂG�����K
�S�b��r ~��Y��u\l�~A(5]�퐡�[]n}Z�qʒ?��
i��`RN������_��i���,��yO��.�����=Y'��9ؕ53�n+sU�^�;��p2(���Ĺ��8�q�sF@����'W�d7;�#dw;U�r��i�Ͻ�erxa>$���9@���yOy>���ߡ�݆S��h^�hx@U����dV�R��H僘V}�t���ⱖ�8Ks���E^��Ԕ,r�7�0���|�W����2��F�������|8o��*��덻"�F���I�Ĺ�P�l�,/��:��S܈z	�̒t�×���\����9�d�5z����Լ;�q3��sť ۵�����8���ŝe��D6,�������|�Pw[��T��o56���khRGr�H4�m>`nJ��G)��`����:�M�;М/lʏ(�RQʻv�@{}�4Gs�9P菇�2:�I�ͨl	㙯G(��4����z��J�j��7X��{h(gF�[C?��8���������Y���![a�%sU�Y*���ʷZvf�oL�c���m����%6]��Ļ�d_ҟ1A����l�x��
'�p��V�KŴI҂#�-�u=���'��f��R�͜�]��6�2��.�;���w��
hFH���5�2����g<}���~x��#v��t[�K���~gR~�U�}/��/>+�}W�4�Y�u�y���5��*�@?�3��P�ZcՙW�`� v#@dn٦����ZԢ���.2�:yq4D�c���2Ax����Q��7P�ag=�Χyu~.�7�a�Q��Ө�]x{S��M�۩� 1�q�+ot?�Y��c��t'-�#������k�]S��
�ͶȬ�N��Mv��s��t�n��R��p<\@^\P��
��������a��������Vk�&��ai�]�H�5���[�f����L�$�� �xb��;���B6? C�r���L�~�hG
�"PZ�<���fo�Q��2�c8�2��D�)��X�����=I��vo^����S(K�[Ăm;09�M�Tr�<*�*�T{�� �|f���&��j^_w�|HY�c�j��Z�l"$t�D���j|@��~� ���'=��r4�b�.A�!��#x��1縦�\3.�#�R"]�����?(g`F�l�w�k��+e�c���olb2�B2	��"�שB��g���B�����$�Yce��|@������,)�\��G�w�zw�X�T��8����'¾8�H�}ac��o���cL^�)��F���|檝Y��r��G�V���ņ�[W-W]kO�.u��:y|<K-7���ty�Tw����`ݟV'ơ2<v=�w��PX��������(�^��q�ޚ�Y�����lRl>s:����Hb�g]3�bsn ��p#��f\zO�N�O�eo�0SH����;H.� �z �ƎeS�E1s"��2�~��e,qi���̞7z�����9/�����W���<,b��4g�	���R��Y7������3~�ц�h?Z�%��b|�m���$�� �����B�d���Dws��ak)�p[1�Mz|�J�Xi��=F\Z��^�.�!.͇��(��gԷ7������̾+8/^�k�q�(����]�U�TZ�S�l���PK����mȼ�$h�'�g����=�`��q*^����N��d����	}�;!���A�U�8ǘ6ǰ�:SY�W�=cf�{�]8i����@ePl*&ȇ��n`�J.vC
2�m0��(�hbcc;����2�?v�%J�i�'Ԏ����Vz��x�3VVl��f��Jn;�[��w�5BQQ���Ѹ�:�t,�~Oz��}
��͘����̀}�sY@�4�Q���$ �ݣ���-�!�1��i�J0bR�^�Ɩu�!u� ��=,s yI��49�"(Ή�ZtU�뫦��"�k�������� İ�A�W���D��_���mݜ0�z�{�9�G���� ������j��gj2�����l�j(�۵��� �P����̹[�܇F[W�.ܻ
��{-]�� .��MO&2D>�5��Z_-��>ӂ�vE���	/��|��"堬�Ƈ�v3��F)E��Q�L���F� dkvr��1A_�) �������'����X��@��p��'Ov���;/�1At=�-U,tk�� p��+��.l���`�"�2Z2֥�h��$�Ǿ%�����=���=�~y�?�̙��������%Ģ��@S���ӛ���>�J̚Ԛ�{f :Y������+�DiP���W���?���AAt���̲��4�C~��C�"�湛���ư����[͉�3�t�_-����ô��~��H�_�$��l�h���20K�A�&n nV%S�{��}6�t����SPTf��<���Z��I����@t�G�H�y��DC�GȬq�jď8���*t��D3�/gfg�i%�n�,��ک�w3G%�n���|([�f���^��9K6�[)����&�F!���\�N���V~x]cq%"3� �ڦ+�H�Ո�x�:#w���B��E,�,PW`��R�����^�᭍�l�X`��S[��'0>=�����f�I�����RĆ���u_Azgٞ��$����{i�[s�7{��17?�|��"����wF�!�������8���
M�W����:So�7Dǫ_�M�&<���eC�˳��lp���X��S~������Ia
�404��|7�1�KXR��TDD����0&�"��(/�X�qQ�Wm��u�!�0�;��
�2	�h8�\�� �lm��0�ww�S08�1XL=�a}U�;�S�뇭��9+���K��+��F^�����˗�{=�:�Lj�
����oЎ��N��z�����$ō�j�;�Vi\�qJdF��"�[����
�� {���EԚ|�[�ž[�	Ӿ.�G��n��KKp��,	~% t]�Ҹ}9i��L��b$��b���m�2|�@fв�v���5ZfJ�}����T�X���u���B.�fl��5�c�3�=\êӃ$!�Ǽ:
�;��T2z�W�~��RZ���{Q���C+��HhUV�jʲ�݄h�s��׋L��W���bh}FC�V2]�I��&�؋�nĨ�o�qpP�Ɋv��%��b��P�mu��Oܙp)�IrKr��SFG�q�[>���t��������0 ��9�����e�J��[�4^�\��0�c.�Q)�hoʥ�?661t����
"���4W���?��3�z�Cxnжp��܍��Q-��_u]����4s��w���10�v��՝<����@y�e�#LW�QgΪ�u����z�J5 )�g�޹���g�*S���I>�Q�N��C_z�3t�5��8}�|f��ጧTVM��=H� [�R�\w�g��_���Bޔ���G=_ג8�E�RZ�@0~�W���&�����~��d�I"<�su��_(sų�Ӿ��w��K��`�b�H$[�N�l*T��f9�͚=K{����
:ss�5�|��8K�r9#:�Z�����y_H�H���Տ��z��6�W��QJ��/`�Aν3F�B6/��� Wj��u�'��t��
���� r�S��MB�+�J������MJ�R��d� ؓȸ�\;{V-B$L�ӳW;?�EQ1s����	~�<Qq2�lrs�����3��3�[���q�,
(�����2Kog�����e�-�ǹ���k������u����;`�ǻ[�(5�c
���D�C���]ͣ$&��
k�8�v��3�u�ϰZ;h_������t{��W��	��H��Sb��q�ga0z?^��A�s8�w�03�ڎ2���ہ1�T�*���*kP��P�
�z�48��.ј���t��*aO��[��H��-�9X4����;aЭ���,�:*�,����T�>��bY�У�GYl�����&�%�ǰ����{c��XU�ږv�9;�9���ip!.�')�֛��s]c7����8g�QU��{7㙆.i�
4q.�P�4JBWV��| S��l����Ϥ�`\��M&�n���i��%MW�7�������>�3{#<��\]�c��M�@�/z}�OҢeg��A�1z�,6�57�V?��C����q�?6��6L�+��N�'VGA�oWj!��Z*HP��S	�$b�2��o|��s�DV=f�9 wBe���8� ��ۜ�í�4&%���~������y���#�>@qډ��Πǲ@XfU�u�ស����YOAR�'å.�11�>��L���0��H�q��U�C'h/���AN��OSO��������dxM����(!�q�I3���2�F����}��=54�[y���{�j�z��C(T���B��~����w��Wed�Ӫ���e"(YA
r�U�]@���xV����6�E��i݂�P���P��B�"�@��Gg`���� .hR��� �a��{�n�|�߂�z�ޑ����◲�;��l]0�=�T(8O���$�u|��J�� .�B��,�[����W*�
�}/ۘVPQ�fmf�8��(b�=�=��I�����\����s��F[P�# z���S6����p�B���������|����dN�x�v�݌eX��J̉�C3�ě79�GG��pm;��e"�����'��[�U8U6�o�;�t=#�}������ �Q�};g4T+N��c4O_��/�:ّD0����/�-��˯6��1<���d)#���[�ck�|����"FJ���
e�3�qͳf����+�VY�Ӆ%GH��g��`�
Q�9�X�ҹ��L&w�"�;�6�P�k�M���P"�{�߽ �0W�	zٝI�|Og?ݍ��h�1��F�>p�@O�5���V�;}:��0o&������){˞�"�.�{���bj�Xe��9/���1w?B�Ez@�NЉ
6^��:�w�!YR
�ߜTf�R�e�+sSVT|3���S�1ʺ�`�nzO_?`<��΃���m6��?�E�}�5�Oz}�{z�-uW���hImV�_]�샇ȝ��ll}O��E5�9�8�g(��G~~A����	�-�(�V)`p����g�JF��{�|�q��|�������� �YUP����yj�޹��4���^�=�u��{���ի�t�[*�^����� #��eru�p����ڞ��\�B?ZY&��e�〤ܧ�t��j�v���Z�$��_��Rq�WO��ߒ �*�����0��*E�K��!��WC{Q	��HO�-hlk]�5T�2���6���x��-��zl:KvkKü&}��c���D��s���C	��F�x��GU"C��P�M�t��8�Ҋ�N0oz���C:��7�?Aw��(qp �R*�8�
��=��{��:�r� ~���n��-�N�5��B	:N5Z�n�O�x���>����
��r�V/����б/�k_�G=N�`�"	��4,>��H��)���pg�K�ᲆ�����nx�@O~��>oί�_\#q�L>{|��kWA�����J>�䅘�V=���r�۵�+8���G��H����.�D;��cJ��i�&
S��>99���WA+��a�cn�ﾢe2��3�BX��&���Ҡ��L�ׯt8��w����� n��.��oh�=ǫӘ�F�$h0V-��+���������(�B��`qYgSh�}�<�����Bۭ%z"���bX=��������d�rL�%��);++fC��������PYM0�g���Ԛ+}����U=c7|IHH`��U-�wUȄGX�>=�8/qm���p��`�����&?U��[�oH?ϝ�h�Kx����uXP�ݛ��fu�f0���/%6��a&1 �C�ۆ��wmb����=��b�۳g�XAg_>h�dP�)W���e<�@�������܇G��S�s�����l���|��ys��f�%��mu [b�^�ŉ:~��i�?�ljk%bz�
j�,�֧�o	�:�֤�O���� 3a��Q��$\M�S$�D��[iXC��7><=����Y1ݭw�hi����Ʋ-ʷ*`�A��;�?xɶ�����8�3�7� K�B��+g�b�҅n6vK�!�<Py�Er��.Z�tg=�u��l�p��(cF479�ea�i��g�|B�<�����������I8<�B ����99�2��5��]�e��.�2��~���r^2BKӨ!��9��g�}|�8_����+]Q� ��9M��"�7���<Ck��t��FS3�j�ߔ������/$��30��x`����D
���<B�Z������V��Ʀ�{N�dC~�x���lgĄ���]P¯���u�E��Z�o�
�
�9��F{.�X��3V�1�׮d��v�eDr����1Ň�Pv�*����߽|T|u6E�_�gS�T�:��bz�(N������ɻ{S����7��-
�0f��y�l\-j��#wE�{�:�G+��;e��E �+Es>����_�䉗�ǿ(P�l	� �j�*�/=7`����o��z�R��S.:�r��Ux���_��`����%�����K	�)0W�w��W�g		GJ�}L��L�I��N� ��<��sf�� �[�R����qʅy�2e�劄F&��Om���eݮEQ���u�@����O���Q_�l�)
�g_����|MDv�to/�8�_�<�A��%8OM6���� i�k{y-��o���@��Z��n�?>;t�yFA4)���;㿛�5�~fa��ipgcj��:2�R?�B�(�Q ����������<=E��6=�B���)'�/ zSS_��e���oy�L6��A��3��Mn6���xD`Jny�'��Q�/g�d)��o���\��+����b�ws�y��H?`��AS.|n0#�NL<���bF��.��U��0��KY�Y�d����&�n���;2�!�r�����0[+4�*t�
+�W���\5�?� �c@+G	�e"�@z�XS}���1bڑ�7��<�-彺<t�9[S��$HyjQo�ɗ�.�x���K�.�>�@�0�����ou�0  �VlQplՙj=X-v.s12SW�Z��!9�!dj����o-@$�����A�=���ܞ���C����nM���p�m��Vg��/ˉ�_��Lp�����!R;Y#�ts�&� ,��m��JluT��AR�]�X�����3���/�	��ζ�P�3H��PeJ�uζ�ӧ�� k�,��	T�@zeL����%�B�Fg�[}"���)5���E���ȵd�� ��tY{�������MO�{(��)��H���C�f@�>���#�/�"�
�h?���"풠�5(,4;��b���Q���?�uI0�9LI�	����rGc��Z�$ ���%�E�S��bM��������=���>2���"45A�J�#J��Z6�\c+�Z�|��^��a6�7�9�Z��߀�zh�]��W�@�O�}����e`x��N�E�,���Hn`�:��.>�ɏm��UY�[7�.e��S&�U�a
l˘q�?b~�{���5�wiy�)��Z��'6���bbM;��^�?��m�{��C��o��K`{�t���$��q���'�o�y�E�Qgi�i���>�a�b7����5_EEf<>�Sлn�=��c�xmԠs�_��xn�Bg�����m��9��Tw����d�t�#����L���o3�(���SHTKds����s��o��n2�N(t4a���y�Rg���(�DAuOϦ��ԯ�l�J(]�@�zYII�T��O�f�"���^:���'H�� �����ҟ:O)W�%��0��J�+���/�"��ᩆ?y����U�(N�L���䤵��]�Ԁ��B�Ϋ�2�QU���N�n����
�CM1�nh�yʯ@LK*%:��w�J?+>8r8;]6��+̉���
],D�+~U�aץ��Tq'(}�2��sΗ��V�����E&�/%���HQ$0��3�2�0E����Z��߹�� Χ?>=���	G�� �^9����@A��T*���<�����[i��N}�ME��������ڋ�H�+����Yq9+�������Qg��7�rP/@B��WP� �K`"�D8��}��j2�'������cx�?G(s�%]��uF�m�߁��CPV�5(���F��4����y�w��Ґ���=�%i�^�Қ?��˨��aa�u��;#�����ө�6l��k_~b��o:���N��2��Kh�8;]!.��kW���<��&K����d��ol��Y������L��ZSb�'��F�2�h�����33)c�����|C��L
�o ]}V�q��M7l�����yk���o�yV�,M��Y�M�\X�4ppĭ;����]��� �m�!��*0����Q_G���a��E"��֕�}wm�����ė�f�X�oF����u�_g.��HLJ�P� 9n&��Omy��RJB�̳��Q����A���Sg{�C��#��A}Ǚ�>M��J(�e]��{�����;N��l�\c$�]��b��c�(��?դd��
��nݣ_?�1y{M)�F�^,��ʂ��K5~Ʀ�	�!���Q��$[+�E�e��x���*��n�	��T}iiJ-A����fg��o���/�N`>Gg�=���ӳ��g,Єfn�ZO~��o�}����? ���z�Зb�+N��Zx��`6ByIYR�?�p�� �h�P�4�/g�m�EJ%�.���<S03f�k�D�OG�q��򱎈���CS��/��xa�]���s"/�;<�<��6���fe�j��#1 �S�II�+�2�9A��z@�X��/yi��4j�p����NB�\��S�D��k��*� l[�߰���Ï`�e<ut�d��{g:<� ��UX;������'.[�I�K˿`���Vg'�ԖWQ�az�=�[\L���3��ou9�n�J��}`�_[vdH�7*���qw��k_�P����IM�{#��L���B�4ہ�˓NLe%^����W�-5������:vw�r�i�yA��.���{7�M�N���~�w�o�
p]������K��P_��|���6=�����s6?,����,ޚӰd����*-c���(rFZ���U���N�����ላP�)���0��!��rCX����1�(%G���g{D�����f�fF� ���F5rbH/Y}{��fcX��j(��x9�03�\��oL�?�g�ȭ��ѹ�ա�*���>����x�ԪE %�sfֲ��|c|�Է�&����HyӈN���>�ۖ㘺Øz��i�~�b"b[@p:3k�K+ ��JT�����wQ-2m�"���g�����9��g��F�G�����V<\�;�ʊ���H����Ր��'9-&\!���8�[�Ft�U0��D�}2�I�bc_�?�%w��7������%�W��!te�����Ý�`�}Tv��@�Kee"讞-�pn���F�q�Ag*��%���T��ѻ�%�z@�nq	%-����'r+�îO����8�X��Z44��7Xc`��ŉl��\��N�{ދ]�w2>1��wW �9����&&��Cx�!*����~�m.��=R `��=\�W*�j�}�c	��22����#&	���")�Fݵ7��� �0D+�������A(�)��"�������t���E���m�9�w,��$�:���#��M��i�y�4g�� �)�x���ra=� .\n���H�brr�]��:U���^.BMr�={��LD�'���֏��~��>���ںH�=�%^?C��U羺�J�J�4��X-o���&�-a�S^�qyG�r� o��U8(9ygz����t��A�<^�o+���~ �h� )�nV�����{z
WcҲI$@\>��&P�r�ZLlxF�w�30� Nr�E0@�Q��8/��3ߨ�_U�6�P}�ʊPO�'�c�$EEl[R�IG�Ԟ��\�G �	�M�0g~������tĒ��	3�4~�]��%T\�\[[BC�SQ�<� ]K��n�)/�
���5l�hT`m�?T�@ ��>�O����q���b'� ��Zv�#n�̌_F6E�H˪�~*x��߽a
�76|����� ���ٙ��+E��0��{==�w�J���B��6uc	o�;~��Y�蓰�ܜPK�nc=eO.8�n㮝��� �j�	�g��61q���S�Q�M޴q��Mx���*�W���. q���V���,��?����xy+�#Cԭ� R�3���ƹ�&'6c����a��Ҡz9َF��,-�����[��6������3u�Q~��Ri��:آL����a�3�D`�w���-���/�es�Os.F�YM�_��`�ژVJjjʮ�;�KX���U�X�y�EYVߨ��ӧ���`��~xϷ�"NGd��r��V;V��eώyf�,?�r�����jθgE�4��60h�ihX�˟Ů�<k��QSC%6P��ڴy����T{;�#�y���J�ӧm@�L�
�P%��h#GU���@C���^���(�+��x3��x F(�|g�D�&�;4�����Ol@�ژY, ���?����3{D�����+�!!F���Cz�m�L�8R�X3�ﱈ�_�'r�K�6N�q)<�efU༢�K��Oҙ P^�˜k����N��g� q�-��7of��Q^��{1���3����huqqs{r'R��T����5Wx��Bs�[8 J	��M������ǁ��Ύ�%���gϘ�n�L���VP~���W�+���U]�;�}=fqW��Q��Z��&���(-���-��"�#d�:[Բ�PR�J��l-?�VOF����t[�"��V�qY݀��D"'s��T۳A�>q}SS8� Gd�o���a�zS��c�D��NSS�Q-QSK��M54H����h(�e����햔:�QK��[�Y���.��Iʞ�rS��HK(-.ݨ���5� +��1eG%&����IK�{:��\]�+�?{uIw)X0��$�|Vt5/osK���+M��sdFq���sע� ��e9����d5��F霼��Rū#T��U����hb�ײӦ�aiU\\���s��C���q?ƿ8���1���-����)滛"=YY��2j��y��"��j�%ݜ.�3�'�4r��� ۝<DG++��gL��\]Ӑ�{��?�x�7�A� Ô��Êv�t�;;\H]��[�^_�������\�w7�ݽ;����I�y�($�8�ˠ��ǎ���Ϙ�q>�+���&�l�:u*W�ԁɅ)�XZ�Gӊ���hb�Y��zcs0�P���G";���8;�Vդ�[��Xpw���:���"]W�9����:a��yOC[Gf 0I�p��3�ᳳ."2ȧ�:Q@���x �'����H��+��&��1W���3L�'`�J�]*jmhx��7K\m���8��ZZ&����XYv�!�g��:�,]D�������C	�\��V��('�:zD��bz�l��j\VցD�DyR-6�jxT��zd�`��,�lm}��^dhh$�k?C�Smh����S���w����/7T�YE�r{*�? �a��:������i�.��z�N�LaF�P�Hg��?XGq����mxex:��%���33��x,�{u�<�R2]qeM�r��z����Q��E�`����"Q�V��4�/_�~��?���
����g�05��o=��ػ|p~ߺj�<�`L�����a_��z��Ƶ�f,��E<�%׿&����>�_$44(ܢ��1�T)��$�Dk4�X�.x$��Еb'|98��4�L'+��ϟ�%&�����$#������#� ϒC�ߟ�Խ(�0�s�r�h��W}�I�3�R{Ȯ��j���OK<b��	�'Z1�.�n�E3������!������|aAƊZ\xCOIT�p}UC?R������o��H����(T��#�m��}�T���i�W��1Pkt�"XMc��~���ʽE_{�*du��T؇��Fk7T׊1�ǖ�L�0}�ç�~��3��b�%{��!�,��yr�$�1����Su�u�U%��v����Y�o���}������*@�!<�jP��R�=���!�;!y���`F�o��նr�f�~=]��>�Y�c%�Q�bK��K�>���.��RD�t9�k�\��{�M4ΞF��<�H~�P鏉��h��k��Ϝ�z^���U���q:*Z\yچ�z�gzh{�C�[����޺�램��� ���i��y��**�����P�Oc�!��q)�{P}��>~��q�ܢ�U	�|��C����Đ&jB����w����.M�0�I|�9��b�[� [�gOk�/N8��p�v���`"�$D���҈�X�П[�Rƌ�ש #�?mja��]�j����@%]���߭�yP�g�3|�]+c�MA�A�ꡖ����iS����`��\�ę=�w�y��؏�*�T�u�Z�����U�ɑ���k��W�=����J��[���󈐀-���m�(�2�Z�x,�r���渹K
3����7�O�s�b�'-E�Yn(��|��_�ǵ�Ja��n��ǵH�i0��kt�JM�����
s����'��8�?[���k��v^��v������;������;������;�_������5	|�a�
���;��؏�[?�~l���E��ߏ���'�~l�����c��֏�[?�~l�����c��֏��/�.{,�����+�n���h�N\=�W�	׋1�1�
��xo&P�\���<TQ&Y�q"Ź/��ގMH��R�;iy��������˿~������N��O�Z�����1fj�]�4�-�+�k���L�a��I��]���n�B��������^�+���m���BߏS��������){]З�U�|�Y����7zz��꼨��Y��=�)�Yk��?}M�jk�a��S)B����s���������tA��*
}%���t�@õ�9�񋰽�,4):3B�*J`���B��e6�A��o6�o����k�.	��D���q}�������>���o��M����.n��+��8r�[�����.�yM���|�C�?<��}�qrq ��7��/�m
}�:n���̌��o�µ���T� C���IP�١\*4�ۥ��4�b���Ŧ�h�>��p�FA�����;ڧ�//]����tH.n����Q�O���E��[4:>�/�}ʇ�����@8��M�Pl��� �4�$������U�]�y�A߬p�ɑ����B�{JEK.�߾������LE	�7%lV7'����τKF�u�߰�y�;�d���z�ף㟣�V*q��/)��I��Z$��צ����C�B�����C���!�_@5���(W��(���v�Y���\��k��Y�i%�hx�r�?���e-V��S�8lv�\^t�W֣���|�.Q���#���@Ay�?v�e���VrBo�	�������YJ����Q~ڠz+Ep���;u%����;ڿI?��B�9q�M�+��4�O�(��ۂ�d�v71�g`�9H\Rcww��t����971��ndd$�C�o��7(+)q��⳱o�I��#��!VI��v%� ��1@����=�"**� d��e��"�ww=�+�]O��@�K�8��^�.P��f9tO�f�7�:W_,j�����C*����q����PY�}ee�%���;��u��e��OPS��0�L��6t�2�!�Ԋ�	�J�eqǑj�`��������M��	fbb�8)@P�p'��\�kI�G�D�8M]��4W�7�u-���� _[��g&*�nD�Z �С�Y��X��ᒀ��9o~$@K��S�FPj�7Pm��_�H��C��\X5�+�{�5�!ǵ1ƸlA`�����̲\TM��h�m�"�g ��`%��*����b��am)Z��ԑU��h;8�-类;��B��uG�T�J�`��1�a���v(��t|���V�'wwu%�(2QQ�	8x��M�]!��G��X�!��̃�ammmVV���Co~���  ��'Z���kӔp�ySllk?ӆ�?U�#᜸�?�`�M�---=�d���eg�/FO��srh�A'�?:�0=M�*��P�]�"� �ꈟ%09���T�R��M$w�|��&����C�$p��E�V�"�˰�K�vF�Z}O(V��ZN�е_ @z��J��<���~<�팘�~wR0d|G��ˍ�I���\�X�w��f`�SR�H�4�ae6iu� `���LNFX�p)B�q��8me�������ɷ}�`àOܭ�Oc����u�;ݎ^P�+{�1r�4����x��R�e=Dˮ��~@� R�;�ӑ�Km���ߎ�y�ǓQs�+�oBrr:2c���gԔ�$=�����-�.� *��/��P��Cm�8�����B���?c3����I��$��B���� T�6k
��Xv�@�P�^M�:m-.*�HPv��}�\Hs�A�ǀR��yH�� ;� ��"PR�R;:/�z�j�#��`o��	L�MR��?��p���S,����.F�r�p "�r�ɣc�b��b��N�-�'��GZ�w�h\T:�Z-�vy���G�V@E����)�wtv2�.1�j=�zn�)�/]����W�ĸ���v/{��2�̓71�����UU���j���l&EEyD�$�=B��� Q���#ge�+P2�1���=�	���Afi�8( �p��0P��%�Rڱt�g&���Ƶ�}TO���B郻��I�'��E8 ����mc8P�:7A��^��n~��ys�m�)Z�|R�yX��sH���K �� �')U:�<L��y��0��yj �C�2����b  K�{3)rEE��9!^8�r���k
gAX���J���f{ĕ_�컀�C}F����&��*�*�Y-�l�*�hY~mHNN>��Zh���#��azT��V`*ճS�h �E��������Ǭ�0Y��� y��׸pv@���U��tP��g:�JKcc#[F����815W]�CՏ��*F��h)����g�T�$��
���Gb�:v0�p`̗��!`�\>�.@����L���[���� <fa�<OL��֦X�q�[@�ٌ��1�Ud������Gd�����Ǘ�&
8n[����EnJ��{v�6���	ǌ2T���A��3ZUV��0>��z���<� .aąs��93:
A��:�D�޻�	�7T,��Mb�\\!vh�|��)��������J�j���R�`�TY�(Dl��\��@Ԋ"�첷V��P5
B ���,.,���1(����Md�fNr/���?��9sf��yfι7�l�w������..uW�Ӛ�Q/Q�����u
�4���yw����:��r&�OS�B�:K ZG�3	LC�c��(A%#�M�T�pG�a߻�fӰ�e{$�~[J$��эw34��'��\2�/�d�OԾޢ;]UXs�x7�j'��-�8a�!�w�}�V�ߕ���?e<;D^a�\汳��> ��j��3��O��`)��}�١�|9
j`��N��)���7��9@�f���`^yY����WhlM�&P��'C�jzw�H}9����w���9(�Jm�#>��&�߹��G�-	�-n�6֖���4=Id8��f�~��c� �u�x�<sΉ<mA�:K��[?ɉV������i�R,��5&���$�DSe�YIKe��1��`��u0�qǿÔ��2�!�q~u1����n�A�xa]�%�Yi���D(3uJ(���_��16�i^,�6��v!8�'�el��$?�)�QHXN"U���DW�#��Í(S0��[wz�����ˣE��d�4��Ӣ
=���O�}R��*�}q��I�o��(T���zZ��)�7���95������w�/ 
||�c�k�J�3���b3���p������R�c�w˥�͡��wi��T�cPo�|���`�zT��vH����x�wO.��n��2�ǒ������\qy���3�W!�m� �Rh����@�]~2eTT����0_*5���nB��[˲;��(p���~� ��c�_W �E*��E��2e�W���ڰ�
)��z�ѥ��̢i����
K&�<���v���nkg�%���\�%~i���B�&&��A�y�D��TŹ��սc�"CD��[�0
B�)O��o*�}U�ݺ������2)4*J��x,&L�qGam��/8�Z�6D�oPk�=��!���<y�$(f� f*z+D�����HR.g\����m� ��<�,0hEzMލ�ք�d��x�rf��4.Z�F~�K�+��H׼�81��]a�oE�v��G6����'L����e�T��>���N&�i�5����6*���h�y��w��#�^����.q6E�Zq�_ډY�݊�y����5�&[�����`-���_Q���k���E��]�Zρj��]��={��5$�S6�d9�o8�ϝ�s��z�m�?��pn%�ХH3뚛�k�<=,��>��R�c�����
=?��DD�{�מ���2p����)��@=^�y-��>ҁ��{��3(�����
[�M��y/�K��j�;P@�"������Ԯ�\�Ө^ZX5�t��"7���V�e�ye�l���?*T`�l�D�3���.R�� '�.T�3������_PK�C�{�Z5�{�H��gKK�W�P=�/�۸�8^������%zz��I�Ĩ��]�($_���8�Z�L�$��c���J����T�[ePA�W�-n����i���m�YMt��I_�@�h荨b��҇p~�ܨS��䘥�U6l����DS��!//��I��d�T�*�z�Qcwp�p'm,���-�I	�5�F�k;���v�Ռ�u�?�ZRS6t@��+��%}K̻��3�+"㙪�S���Kz� uv����A�l2�q�בV��<��dk��z9L�Z�
'�n�R���b�4�w� 1)��rp����gz=�?IzO�f�]o޼9XS]=C�`��=���C�1��B1M���׹��5\���'_w�b]o���I~5j�t׫��P��u�\ۼM��(USv�p��p��P:���{E�w�׉�r,�78<�y���i
����Q�\��&��+��`�IB�u�hx+���_�����eb9���'�QķG��wqr?cD��Hz>%:5�`�0���ҝ{�t}U�D~��7����	�gɦf*ԸK��Hw� ������_�>gK���^3a�u3v�,p�h'�x��J�H��aN���s���������lIp����)֥�pmF�E�����$4_Y�Xߒ���Ιk�Ԗ^?�e��`5[m�$��)ƊL�"�Ҁ�����89�e�y���X`kY
_>s�����'�Η�c��}6�}b� iU"�Rm¥�Ӈ7�Z��N��}�.ni�E.����[�,;�ߍ��]��<�c9�!�Y)��8�Y����$�h������H��K�4}iU�Y��@�tॏ��Y�9/�8l�x�m2�]���Q'0��V��?�1μ�>�A�;�dȰ,��H�i�ĸ�E��^l��
d����o=^��-�x��	n�O"�������M�F�6v籃�mR����(����!�W�T-f�3㵼��bK����))����E��%دcc	Z<uh5��"��\��s�=	<.��J�������C��į�Q�L���c�!���B��jL�w�<L������X�$��5+It*�����'��LU��� �P�4�P��T�"��������q��I��h�8ހ��c�C?Ț8P�
�$b�2���<�V��S:8z�'�u�H�l�_X�o_�4���?Y���{��s��7�gXֿ�b���{YE���߮NO[Z}��__��u��k�������W�t��/�}~�r=�.�L�c�qo+?�*è�Vm�ќ"���Qmc���_+@V���]O�
7��}���i��ɓ'�$�i�:EfO�BG�y5'�[���wg�tΘ8~�b�=.ەi�~X�g
�K�a<��d���p����P��WۮA��3���jhd[�#t��-;������{�"��[_<��\~��օ*eKa>�$�$"�G�)NH(8<?M�H>����4�./��H=���7���t�yc�#!hU�i�����[�N4?�w��؅n'zӷ��v�-;Ў�AP�w=7�KGy�)�����x����H.WhAƪ�(~����F	b�ɅB��O�#J^Ң�$���P��A�nQ�-�����"��ϧ۴���~���7�\S�Qk���ؒ��F[H�O�[�`w��fO��zG{ޥa�)�l|��Q�l5�竅D4�"
�{��ʤ��?p��W�,Y�`�<��1����\nQc�!ˍ�z57��-Mt�_O|w��rc�Н����"�kɳ8��������(T�⤶ƢQ?O�٤1[�}1��9b������L�|����������}~V���Jr��+[����-Q�J�vg%:i�#1cTQw1F����0��� gWȒ�---}iJB�_�mHN6fv>���gXT�co�=٩BgM�=�Bg������Z��l�AvM�y�ۤVG��p�� 2��w�L)'�b!q��J9�� /�]�h �y��
�z˥�ÞQg�ImO�Ԭ*QC��}:O�(A�+0��������M�J�f.�!L����O�0�ߝ�ȑ����*<����AuuujP�9X�^ÞQ�Gb=���h4����>cSJoa�S�2���B�z˪"�������lkW���6(�V��0�w�z�č|�ԙ�o�O':��)b6���8�F���-8L$��6ZV��SF��@Ss؇;d�>|�pgHȈ^�*��3��*���ǎ��Jf�������J���s">��(l�Bh��_�t���C��)$x�Q/�^7٤��m{�YfW����:v�<��==B؈���|�Z��|�L��,-3�B�p]DP.*�kw;���s �MzxyQ7�Т�Q(�F^�d�����k&�=�e���\[�����k���]ޕP��N��W�������G�[����j��A���+E��|���~X�@��8���L7�����ۥ0b�
��w����"Cm�w7T�I|~I��gݻ�Oij�Dyo�E��?�5�)�h>��kd2�������i�iɻ�H�xy�����s��
GmqQ�o@ na��� �L���_��u\xO��ΓJ,���y�u_����5f:��5nٝ�b��'!B�Pa4Al[CA [�s�l��GfĮR>j��(�0S�]͊E��ڥ >1-
�יe
�?5�w�fGp�ߨgv�It�%�,Up�����B#-�<t��s��?>o�w2g�H��82�/��v�^�E�Hff��$uá�D!O�R
٨�#���dN�	�yCh���a�}����F��J�1�F���y��Z�p��I�����W��[���۲��݇��B2�<#P�w���O���ų^!�v5F	��)�1���ʸĜ��ڀ��;�Mir�Z<1����������s��c����ξ��J���<(z�B��)M�1d�k��u��������I�tY��޼��?��#�>&�`^��"�����+dwhF��{�5(�-���P��{ o�II�ƶb� n�N�-�R7�����N�vVjʶ3P��L�(�Rw7B�@��G,�R��J��T�vR^ug���ѣ� ٜ��Go�Ȣ�޻w�Y�;��MwJ��4�b���No-O�wk�S�G�9����9�L�:/
s!���w�.�~Se�hNg~�)>�ȂL|�Ν;��z�6
�)��%��f5OA�S'7>��QFB�E���4.��aN�?q��?7��tM=� ����V/�	z��"~n~Zk
E0���@��R��F�w(Jk�����J�MP������)%S���i_�Oi#�`��	�2<��n��^���0ϙK_î/��zK�WG�2)
��C�ū#oƐ2G���3�����������\!�+A��S�%'��L).�ް�s[��nS:2<8:[�3�Lff �0�ܲ�����F�w83�u ܘ�%����Bn��u���Nl�
6Q*�I�n�r�װ��ԝ^�P��bD�R��?��s����� �`��@8|�[���(�LE֯3CGG��sFW��8��fܺ�Z1��}�@]� bX���G�{	s����2����K�9�(��F���{z��$x9�A�6�T��+n^�}���g4��9�k���Z	6�:���DR����{�i�&�,�Ǯ������|f�)�������J��k���v������hcJ/� ����:@ �qM6��" (Fg�X�{x=�ŏX�v9��
�b?S��� �L���H6�a2A@�,�&�b#��
)kZ���!r:�9���l^���j����H�#�Ϗ��n*�P�u�'��J&gj�������^	[C]��X ��|��<U&����D\s6���~M�dB���#�}ɑ%eն���4�6%Z��0џ)MR�?/��[E�*��O@/�k|�%��s)LW&)�Zka�ZY��j(�] �;qK�?G�l�k�!cѫ_���5���<�q5�)s���d�\��=��-�1��]MԼ��Q��\}�5x����P�&�υ�VO|�_N.��_'1�'?���X��iS~Dx�tt�b>� ����Eɕ-C��1JO}ww���aP�5Bé.]��z��l;;b��n`샱�7�֧��G=#�����A�Uٙ�oĝ��G�'&֢L|����Os��*�W��v[�:S[?���N݁����v54\�)T��ׄ)�������BC�@�����b�0����=SA��h/D��Ľ��Ə+�M�i���9����[&v��}x�#ۈ�ϙ/4�(hx!� GK�^�,��m��0�.��OtvvN�b�/�8%����]��,Gi������@_^�v"��555�j�N&%K�%_�O�$j����qI�R۞��Vc��d.��R�;(��i&%	�o���q��IwB43�Y-��MgFa	�g����N�9�	���$�a��
�F6sU�=�SZ�Ty�=���<�p�I~i�o{�n~"��P"JKk�t�`�EI�C����Z?��� _���?F����@F|��-��"�\'��%m����9��ߺu+��0��oi
�6B��_M�I $������3�~
A|rg�7mU�1~�����0\��$	�n�on��s���7 �����f�
ןFk�0��RB�pB-�٘āOıwRO	��P��%�%Vp���ɆҨ��ɅR��Br�^K�Fs���-�w׎�wS�;��-���4�73��)n�LOq�KS|�mo��#��"��%$aL�1>/J��k�����z䓡[G'����y���3�/����h���_-n�ĴM�9�52"�+�/���e�i�0G}[Pw���5iiD5v�(����p�h;G�4�o��rVH^Ւ�$X𲡸4!9��S�����i?�J>�`%�x�L\�:u���qS-Ε���m����>l�����Z�Qw2�����Y�a�"}��2Hm)��n_��If�C>m|-N @�! ��Yi�1o�[3)'���6�Ό���H�풉C��bn��(�S�l�6��ajL?�dS���s)9�m|�Mu�|��w�K;pQ,'I�=�ԩ!c܀���x���+[b�힦E k�@��Χ*�"�N�����3�� ls�dq~�o�U"�v<���z����e��L[u)��
�4骵�:�;sq�VNS���ýGz�e`��uF+;R��?inn����÷�l��M���JNA�i��Q����?��>5�y	?0Ց9,5���լc��fz���WEE�qS]����:�+��Bф��&YB��q��PU{�{�^o&k/���.�l	�͊��y���\�5#�$#h���a�?B���'��&�����Cjb���s
��7�=䌨�A"
 B�E[�Rq���l�N(�Ĕ�B�dh���S/<�Gaů��v�&�&p�t��"��N����fH/��	�R��g��<c��1��0DކA�̉��c�|�8����Y;8�ػw�I�w��Wf���5P!b�f�۽�L�V���B>o�O �lV��.�{kJUn�SL��>�C(8�@K�M����K枕h��-C���XE褛?�9k--[������b'��L YO����|K�р�C;%��$���$`�v5嚸z8u�A�Mm��{���=�nu�'�D�&%>`���J�����ԏ�;*��|Α�,6�$H��S4��{4iۤV[���	pxlY����|�xj�K���+��3ձ�W|�x����d+��r�gX��ˆ��a���/l�F���|�B���#�P�Bv}�p�����-O���[Ba�*;��0`��=���7�ŷRU�z�z��I��s
�W~:6yv��[0kͣr[��6�-9"o�0�z���:��G#���T[B�*��#�SZ>Y����s���K�b&�춃�Ozc�C?��N�h�pܫ��0rēA��a���6~ˌ�r�Ġ�;��GIc�4��Rq$��#B	z�K�J�^����
�d^�d��ifl��d�L=��tBXۨ����ͭҁ��Q	q� �J�u�]�B�kN����,rP��[�����I�O�h���M��`��/ ^>���֒0=H�bQ*p�]�-x�f�,�+�®F����dj�D��3�v������π�+��Y�=�{�����D�3=�5��B&�\Q�	�>��$ޮd�O�J2�b��iK�o�,�N��e�}�W�)7W���g����)��׵���kB�4f�x���.���$'_��Ѳ�^�{um�y}�:�J���F�P=hM/*�CS�S�|}��1,��+��m�"Ɂl�×�@�mL1@[&xI�I:O��n{zE�Y}C]�9��j�������li�7/؈�?a��[��=X��G�)t�*����#$J>�"��/هz�C�����.y���7�=]�3�ض�\i�W߫B:Ŷ� 5��8�oyb�l�7T6YY�[#��_Lɲ�wa���1#��~�z4��#k�/�B�%�Λ������P@�`:��sێ���9�U�h-��
�f*��s���PX�Z?��P����ɌMh��$�K.�����'��bz�zrO0/ �]�vͮ�g8H���b-�#h�˩�P<�dسK7w/���J���U��!���+kb?���\�$"h�h
)�.{��9_�^8��K����9w�x}�����O���̓�-�P�7��}Y6��V�6��7�~��w�p��`�Q�<9��IĤ��$�PW~��ݯ
�g�G�>���H�ܑ�hg
~�+�k��2�&���[�6��_a�ap��S[':n|>�M�-oFۙ��"Uf	j�WB�8�cJ�L����kZ3��1��A2�2�s�W� �� 6�z�fiE�͉��e��,�#_a����Ȏh4�N����ѣ��e�T���%�=�0�ҕzK�4,V��N���)�b+��D�W>^�ũ	ƪ����xH��	
n,���xw&Q��l�B�F#��^���-P�O��oM��.�+�ܕi�.R�I؃�t�;�%�$Bu�����YR�^�2�О���@wz���!��<{�<v��t������.n
��G
��^r��cK�ÅE0-�	����Q��Q���i_vm�\��0z<�����9��&`�{Xe/SSSup�u��XA�%�ʕ.{4��e�)���eo�ī2���{�ؾ�e=D���)�	M�zܡl�[U�.ǀ	^=�T�|� �eS
�s�@��	�1�N��ìq�:��-Abc�z#�jv�������y~E;!�_Dl�S'a__��WS]=U���\������hkkc�Ǒ����d�Fë�]�H�+��>|X�Qei�0�����M�Q #S,�m�YV�n�,��Fq�[�O�5ڃ-�k��zȩ���y���^��:Z[@��wߔ/_�ͫ��O�շQ�c�ՓwI�yC�ȼB>#�w�<�传�w��)j�ͻ-����\���u��B���������P��W���R��F���?��7Ae�h�����%}p�ZM�Pi�Sւa���k8, ��z��*K���Hl�-1F����Ta������*���-`�y�M�x���vÅ����n�\y�'�ƿ�fa?^�~����]=��d*���rb�k&8�W2܁>gsK�L�y(&ѩ0��6����x�O^���d�t@�s<���1�5BuY��E�q)�k��=d�z�F(0�:
�I���@'?逦��9qѣW����y��m�+�H��)�,f�6	fv�S�Q��ᐢ�G���;�r���[4(^����I��9N�3|���f�1���+�1^l��[�W_U����vZ��-.NW�{%Wzi-k��+����J�&W�������w�)}{c���7_ٝ]�W��{��O|��-��EM����}�hZ[�Z�� ��s����t�\.׮�[2ͤ��s�{kϑ�iji��`�\B��#��o^Q�W�/W��)��y�!�(��H�F�Pb��MK7g/�	�/�a�pϓ'Oҁ�����ȣ!r��h����;{P}���ȘD��s����p���	}�;SzX�M6)n���É�NY$0�Rm�b�w�K��U.�.�����e���?c�|P͔�Xwi``������e�
bŃ��-�Z����@)�Ng�2���:����x"f���h�$�Ň(�k���ů�n�['�����Ǐ��kɄ�+T3�&A�>'�"}�`�̾�q�
3��2J9�s�]���cW4O�O�n��_��;��e"�gZw%i���Dۈ����I�j��"�Gݻܐ�esYD�K��| R�%�vQ�����Oâ���l��}7��?��G��O�v"� ���2�HF���ħnj��r�Dۇ�Qq�8�b����O3���;���԰%���,����LOK3��e���a����m�ήtw�qLF��2����C^O2)9H��y:>�p�L��dq;Հ��,�K��ˏ
�m�%!�+CE���)�\l���7�K�d���%IhMJ��2��$nn��+/�t�nS�D�	��}��>*�VBIfWc�m��B�y�l�}��~�ŒU��V�/V3�S�-���� F,'��+z�KK&F�B�m�<R�dxܺ'��(��"lD�o�*�qb|���
���hk��0�]��Y��`K��ml�#��Oe�L ��Ni� 2��/���ܼ��ſS�L���Ȇ��
���6�5�N�!kS������r[�*Q'�t���Z{?�5��R�{Xx�I~n>��gI�U���s�2t+�q�J�}n��Lt%F�P迣�1t����-+%����<�y��$x��0i���GK��a�l�_���WX�S�Mg[�`���i�]nJ�Y+ Ch%gѻ�D���C�&n��m��^.7������G�Oa`�[H�χ��vNR7��So�g�����*�l�ӣu��q/�̸� #�Y��{� �ߡ�7��ٴ��,�Ƒ�
gt�o@w�
&,Iu1�w���l��nZ�2_��A�"�!�|�:|>�FZ�IO��Z�~�?N��`�D�5֎�9�k1[��(*�>��/u��z�@+����Q���n}�h���Vd/ɢ�un�S�+����]E�q��k��a�k����bE-c�>L�:���t5;�:���^�w��<O�+�% ��Vd�c��7#}Q���R�Q5���o�BI�s�͔�!�v��ck"�1�-�v�q̬lɟ)���U��)�8�t���Üv�.��	~���s�4�[(����Ȳ;��t`DV֤�NMN1`�Og� gvF)=5UmW��)�՘��v����}w�Kj�
�x�tt<�r���Vt��	�Tb�&)su�<���D{���K�F0�"/)9�|^�	��2�f"��b��K�y�F��~|�~Qs��3tJw�z2�1E"Ga�V�/:J��PJd!�'��#E,��hG��!�~�Q�;������ %=8��\�%����*��VI�WVV��e�b*&	���շzJ�qK���Gijj.?�@�M��UM�mj�T\�d�[6�@���u3��"B�ڤ��)))I�J���%�Pe����=��:�g:�%x��w�����
�������ȓ(#���p���%
/5V����B�ק�R<y�^:
x�^�^���I�m�=[F]���֚{�3�	h��Sj
�.�*����)�0�XZB�;:��W��;���FԞj��6Z�6�|�}A�É��e��>�a�ǁ�����c�y�6�r{�n�ڥ-�)MR�E�C7��bF렶�𒪓�No�7^P��_�9#�!�~������Os}Z�k��v�� ����_�񸮮�!đ(/�o��Rw���WD�\G �����(�{�����[f�~/��^i�Mu-MMW���朲޲j��c�)�i� ���N>/����m��U��f�1�'�$j�K�4q�*c��`��-{�9I�I��ʀ R��O�}*�����KU�լ�lY���D�~OX�㟢�x�,--���s���~�U�kA��L�7C
��c{m�i~�w��Cn!)r	�8��gϞe��>����b9��r�,�Zc�Q�̶�/�Z�������﬑XV	3Y;��ބ\`�)�iRRC,x��S�w�1If�P Ly�3| ����@n/������xe���)�>���ݭ�]Ky��ƺ�ӧ�Y vz�W���
	9A�P#�A�Ѓ9@��{h���-tڱ��}�,����&n�ٚ�zrp1�����z_Z�U%R����I�ۏI<����]���LN�eItU�1;����ӧ7/@���%�I�}Nh&����hIͰ�*���?�5O\`h;�	�6����>��C���_p����H����*=���Oڢ�=\h5�x��	�?�*Lw�J���A����"�ҳ��һ��W�T�tu��s��/�<�����7�dK��d^����x��{�t�$�^J)Z��"2eK���Iyâv���T��G�����w�"��
ɥp�r DiG%[x���	��O�~*�％��qhѐ�~�wL#I&6�I��D��H�֯�Z��^����+>��wEid��̖���u��o�V_I�Ç�u-��'��.x�J\�?$3m$'�c#��W ����=�'3����99����t���PM�s�|�l$��͆-il�0�r/̖�ʲ*��yVs7"��^��4����YjH���8 ��!KEa�P�g>/��oP/�QeQ��+�}*���k#兑�,�����[�v3�m��r�����z��t���ׯ-�΢_�=�)�*9�>ګA�y��U����2���R�S�̄R�6�Bq��/q�94�ï�,�����2�ZEC�1,�ܧ�*�RgSJ�EaN!�W9�=i_�H@��tG�ֻ%Le����J�`o?��h9QJ�`N	�i^ҝ�J�s'�x��63���>v�סd����GF���'KD!EN1��:A�9e�e,-X�vr'��`�yqwh���N��tzN��v��1G�+Q'6H�Z��\ûh�ik}]�������*�Ϋ�o�B�v�B��sꀗ%L��I�\h�*���ak��Xc� J-̮�dM@�*�}��N�^e|�d�Z-,,d�_�Η,�0��:Ρ�	u����T�U�,�ws\���Ȩ���5>�D�Ә&D%ǒ(Y���dVٵs���wĹ���)
-"ϓ��Y	&�jw��@�>��Py��%$��]�~ɕ-A��݌�ɆHo�����.ج�!�zD�����Ѕ����{}p�y��ڝX��N7�����5����<�/٩G�M��dD�K�������/�|a=x�z>,A��l����g2י���ٳb��-��lTH���SKK�#�J�frV��\[H�D��MU�!i��nj��>[>�LM��Ԇ*�Ϲ*[��|�ߊ����{�����0_J��/����T[ufƆy�� \���3L`G�a�o��)Yr�oPt�`��=�r,0��ݳX��%g0.8>�}(�����n���z9/99M(L2)!��rU}yP��+�.i3f%'xI�T@�ܷ�0xP:K9L��9���ٵ�2�S��䔴rGw���*�cդiH.�>���~�.* ��H�FtI�����p�KLyN2p>'t�C�tl��j����z���NU��ʽk���G:�y�ƭd�B��K�C�� +}e�Q~FqbL\�]J��Y=�)���uq��9���4���eW=QDV2��jM۬-���cc���I�3�5	C���Y��S����ROi�Ye���ߌD�1���H��}"u�8���<�L�*)'3��(������ u��������ڎ�`�r��kkk��� �J�~�Q�qdA�x-�ɰ��:��n!MT܁c���������wB}�k�)Bs"�͂���^����ID�$Ok\�l^R�&;@���Ν5`�	�RR/����ͫ�F@Ѥ)��Iy�~e��*��%���3lQ�ѴvW�''�g57c{��)�7���83q-�l0�Q��F3�ڇ����Oi��p婴����swϴ���d�>/��Z��ݘ��ԡ#�1/�r`W��:2�:��ws�-�����Ɇ��X����[�D�Z��*�0����y�Gp�+�4��$=�)���~�����$B�3�eH�B������0Ԝ�M��B��k2�$�g�^fW!�Q�	>S��m���W�W� ��$>������>hb(O0�T%��%��=�3�����Ɛ�hC]Yh`�������4�)��|���m��Ii����E���yk��U���Y��H���=<ğ������yb��B�B�y�-�B�ZF��O~V��Q������*!'�w�} Q��	ޑ�1w��jFX3ԙ�İ�eG>��χ����C>ݝ	�E7�zDT�u��3[�H�b>R�
��1w�¶?Z�n���#��C��v���N^#���X�pA����:{�厴��6.IB��$:����<�L�Z6�'��i\B�K�JB]�,�jL�8|N56�@A���Ax����=��s݇��cS���k;��6YY��Z ��������0-Z�og��Cq7��k�Uq(�W�nT2f���۽���̮,����6�m؝�F�r�=�T���aNJlݟ�`H5��*�s�y��h(�F�Q���PP@����C?��MOi�۾����u���f�c[Yf.�5�A������G��<�~��߹��(��Ogs�sds555��Si4����M��i"��6)M��(����? a��0�lo����vt����|`6-�R����*TT��,h��C�v@��1�Iku&w�|�ip((�&��)t0��$�k�%���la�k�Î��K�2�W{�)&R=|e.xρc�e#�===��(k��u��o^(������tP����g||�?�kqT�}ܒ��m��Vp�����TQ�T_''�+g5�[�3Y�{����E�_�*cRr�&����%�r�ȧւ�I�p:���\��x?��Ǘ���u��yG��)~�牀y��<z,7��]W�����5"}|W���ں�-��*��[8�����5�3¿�;A1j<�ѱ��E����i>��k�tP�!�ʀ�.���Ӷ����������	M�
1ëX_��ЗDlkC�V�rZkQ����D���'���ebL_����7_oY5��܆���4��4<���� �Y��s:���]�K������k��o�U�Yv4B��ni��յ�1ޯs9�)%31<6b��&�.A�}�%i4����W�2M�NF��P��台�X�l�jV%<`�Ѡ?���<��s�Zn���������~�� ]�{1��hZjj�Ld:�٢��-!�����������|��BE2����3Sa:�!�z�z8�³5�E,��+l:���#H=:�IkzVe�福��x
���$Q�r|55�;��
�Hm�x�q���K��k̝�?GL�f��>w)?��95c٢E�9-�^6/BM}���e��w�Io��~~>��\M���KC\�٧n��8�=����e#������"��y�17 ?�_�~���5{y0p�'�4��q4$P�8�T�ꄃ�z�S�>���_C�p�t���t�UL�M<�3�Y�����.7�sFX_��liiI:1vj�P�`i�wb�1��<��kZ��C�w�eU��R|�Ӈnc�<A7�%>y�)��n�XOybH�����;+�j ��!��VA�jYN�����'>�\�s����Pt�c�6Ӣ�Xȷ��w{�\(�/�c\;(c������ҒٕZ,��;�[�0��G�%��D����OvgگǗw��*�~�)��p�_��[�C��*@&4��ݧ�A'�sbbb����k�ل�ߣ�`��i�.BhD|��h���#,�Ǝp�ִxO277_>�e��EY�#kO�������M��u�bSB&6�'#���R���TIg,[�Ty��ah|g?�2��HGG|�_�	���R|������ii�Ȳu8��昁ǂ��d5�8a/��!��8vj\�f�(l\mB/\��D�pb h��}�FwH�0��i���I������,�i�6!'�=_6dj^9��>D��YNn��<IO�P�@�d�ڬv쀎P3f��w�(p��jw��V���� �GֶۓN�8��Z��
�N�;��sxJ��'k%���C!k
�iI<�ÿ8��
8�n�R��ͫ��w���&%����%�˿7A�Pv�14�����/�{����IY�m[��U:�z�����7���w1Wk�¬�*,v�W�ε́g�.T8F}}�3%�~�u�p�x�������C���Z�̼��;�����㠾�Gy�95����/;��[��������~�e�n]@��4�j�������/�yٵ����y��w�ZeK�6��UP�?t�/޾;�MD"m�0'Z�~�e����T}����.�Y�Ź`kF)Xm��m��i]��+&q@��9�e'h+������u���RO�0��u��.W,`�^4z7fgg�U��U�h�=���7>�	�`%>�d�ȝ��3Fq3�M��Í��N��6�1�*������hS��-�;=.B��;�ᒖ���{��~�Ȱ���3��Uf�q�ƫ�� ���`�4%	���]����3)QB9U3�����E��U�����/��̄2�	K�k^�����J�^v��4v-`�h�U*��^i���������ސ��O�mS�7i���Zң2�!�ʀ�>�h6��XD����6��a=�m[�M��+��o�{��jq6�d�͓~���A�f�k���\Xi�3p�!����ͻ#lZ;w�nu_?y��4G��t��X���F��3�.=۟}���V�����������*��*S_%�N#�}�����b�椇�!b�:>X$�]n��BՋ]���O��j��Q�K��c�M�zt0�T�l$Ҧ5��u�[���6f���G���ܒg�yq~SOK����.J�����z�P�F�rS��G_Jtj���`�d�����=@�0��wcn�8����`�����������?�e������%��x�J�q}�����\�2���k�x5�����=zT	�vqfu:*e0���U�Ɛ�������$�V�msO���	'q��1�L�Y��q��98�σ�jD����.�\�>m]�N(�+JF� �ռ�|�&5�w�ɘ��$O $Xp�tA��]�9�y	�(}7��t���eqkC٬B�e��i;��;�f����O���'pDy���=�ڷz{{�U�8�1+�· |d�`Ct
;�OdV7��"D���\z��Q�"ufgq��8�;�sW����{%��;AxYz�n�D�hl'��lݠ|~vC�U�7*�N�]��a�>�	***�?;����^���8�C�|���q���� zm���D�pH�\ߣ���.u�Cv諎��`ȓ�ޏ!3�޸�C׼��@��^oe��W1��(�,�ruu���ه./{u�$rF�H�(��A�p�?2�ќa�xJ��$"D�X\��S�|E䩈�w��[���骯rA����}��T����	c���.g5'\���ާ��
MTO7���G��S{�1����<|�O�l����
Kޫ�k�%QWQ��?������z��6_���6Z��f����^Wm�.��ϸ$�0�W�W0�L��,����2��U��M7 ���0���ᶝ���(������#�~c���w#��N-��t�B)��>zl��ߦdV+|�	 �i,�f<8���16���in�4@�ر�o�x?�95���-�	�f��9F�o������r�����94�O����<Y��x���O���-2�s�DdeR�n~j3����3�gc������4�䬉z��I�Y�ٍ���+ �TU&�s�H�=�L�\k��C-�u	(ƻ�g׬vB֮�>����O^UrH����ga;����G!��5K�S���Ts\����ɘ�\:j|>{U	�����o��i���'�]7p�X����x1��}��DoFd6>�"�:��Ym��c��gli=�dA7zbSp�~b�@�?�[����#��A#l��;�c�)
����xP��7����������z�֟#��h��	�:8�zn�����D� зy1�{�ٯp#g,��G�ؙ5����>���,��������ɘq����5�\n���s?K�V����$�1�7�YѰ�	x��`Z���s`\~�J��
~��e��_<ϊ�P�pD��L��^���7:�}6�Ψ�ǐ2\koCX�G��3��q�)��<H�S�F�ӈ"�0�K���K�
g�F~�k��~AO��?�Ҍ��3	q�Ol�I�9&�E��zzf,�1ow������Tvz���|�Ljc_�ZQ�Uy��1B�y ��Ŗ����/�G�u�� -�<�ƿ���
�h�$hث�G�Z�p$��{F���f߂�۪���-��?�G �+[R4�ŀ�u�vw���
Cz��J����Z�|M�����6sA�����1��c8�~�ͬv�$��,�d�1�:�N��Ł�݉՟� ��Km�n�<���  �MA�jL(��:�kٯ3�`Q�}�$豵U�t0�rf!��g]��hn�]���e�^^�k0Fi��}�km|jf�23ҟ�R���FC=��3�V-C�+R"2@�� b�Y�����j��]}8n=����ZSX�k��[�� <�-^�������C�;�7��hGe������2t4vJ�{�l͂�-E�:%���ڬ�˙��� �܋�˔�}J��.����?u�do�������K�@9g�����c[
wuqY��Đ�y~}�������p��Q�;��g�%��w2+>�����ID����&m�?��\q������\2�?�e?����ask�����7}�q|���wà��N��C�l��683����C�cf��R;�p��~�
%ج��+*b*�Иd&[���{�p������|ļ��`�TYc�}����/[veuM���`?��K��s�7�﷏�.8��ӳ!"ݣ�C�ZV�Ǔ�R5P�߯�C��׎��rvn���}9�.��xJ�ec��
�֔�ŀ�]�n��P
��ql�Ū�� /w#^%6)h߅���fm�;+�,�� 1c죌ǻ�Cٯ�A&����g?����@��6_��v�7��vt.���k�y-���L$���%	Z�;�4�/=�(=���^�j:S�I\phX�}%���%��5��r�~��� PK   �}rZ"1^F�� Ho /   images/a027fa6b-1779-4bc7-b1bd-261c8096f986.png켇ST��><d��deYI�I�TT$G�QVQ�	JD$�` �"�� #��!3��ׇ���?�z��*kk�;��sN���������T��e��`0��gN��`�
1��m��\��n��v�3�1����GK=]��^��.���]ܮ8]ø��	[�Y;�_q�&l�d��e�`��UO��s1�%jKq�y�<"����j^O̡�#�Lv����cI]�hz�}>ʹ�S�E [�P`���m֛�fZS�h2������
ϯeg�?���0������O��ӟO>����ӟO>����ӟO>����ӟO>����ӟO�?��ϳ��==�컺h�p�qW��7����6��P���z��E��[o}���MԳg#�2�F��:dk+k����6�K��'��jY����8���$�+��=6��Wf���1���x����>�u��z���n[��|���?_���ϗ����/�|��͗+�j��)F��������:����e�N�
�gV=g�%�6RIv�����h'�⏑��P����!�c
�)�}�ْ��n(8T,�	�PJ�I��������K�.I�y-��K�/�9ƚ��g��9�)""��K-��#��Q^�����:��վt��xW�Pɷ�o129�~e�5��>^��3j6��G��T�}���hM�14����bbbW��3mF�����Ռ�����.e�����f]f�r�˯}y�4��n�[z��6�g�I&� ��o,I5�8רR�����<��[o��E�Vٸ*!;{&��0��޳}6&&&��X�a��\�f�ǁ��,�%�����)����$���|�y��_�=������U'�I��c�S87���^��*���l&���6��uS2�>���M./�W .J��S�����V�Af��k<���'=��}�=�����<n���*�.�O�fp��M֬IƮ���4��_z�E�7b�/�}K\'�����c}�Glb}:;��U_�,��;\���a�-b��`�����pFYCCCL\�ڱ+���^	)ߣ%�tUv�E��ȶ;���Cʍֶ�j~���{��z�5WRB�p$��n��=�,�U�o��_ǳ4�%�e�t�Y��G�O�	eR2��(�U����/|���W��Kbܺ�YS�V�Mu��Gk������Y��;s�㵷c݀u�n�);�i<�sk I�/_������\3�T�_��m�;�?��!77�.r����O��z<�,��.�N�S�![X*�����v�\\]���4Oܰ�	m�R�Ӕ��g��c[�ߺ�A��Ƕ�~�Y5f�uO��k�ۣ��2�jk{{͡��'`^��2`�5�0�KF":���x�hlDO����6���doYB^�xH�"c��I΄�%��%�����L�3��+|}*��0�n�1A%t���;�<��;�m��XSI�Q��l������*�u�0\��}�������7��Ct5����dV>��V�v���o{{����#!5<~����,�x��|��cg�x�xz��g�M�L�c�%.Lt�d�u�#�9Q�Otw%�ysx�z�r�sw��k����v��1#�{�h��'���N?k�f�K �!�����Ds�V�!����!w|�9k�M�v�;�!W>޹�ݽ5�`�mmO��,z�&��Vx;;�N9n��ٷ���� ֹ!�u�i�b;���W4�h���9Z�;g��k����� Ƞ����n���ٯ��E�?�O����[�-]M'�]Cq�Аmbb±킅2�wk�1331#��fS�����n�e���!�Gx܃�Etuwu����{�7�2x�������e�7�>�����R� 5ss�^�"4���N[��9].gki���s��{%�b�X������C>Ȅ?�c2��LT���u�7�QQQ�t��'�\�9H�Ӟa�6�J�֫lޔ��a1ſ~�Bp�ƤL�w����=�%�T)Ӥ�luqڱz��)��$a.`%��ӧ{�]n�N���@T��.R��X�������=�v�ȋ��H&������Dns��V�IB��/�,���x��Xuc�ó/�D�����I�/h��ʻ+͖f�\F�\j_��\g������yu�0���/i_��ɝݳ�� qe2�̋@�tgr�zǞ�l�'vpJ���2�(��=Ǯ�]5�7�����\�ۜ��E�`H�pk4�����>7�,�U�-t:�k�«���W�sq<��
�z���f,�����Gv�1�"gmoJ��ۤ���X���I�����RY�UY��E�<��S���"����{fՇ0iJ�#q�g.��r׿�؛���.7^j6�,����gM���e[?b�$���|�Mg��X���i,���Y��e��� ��;�o]���E�BLR���*d��6��ʲmz��U�f�B�����;;{�uf�鐍ut��S�i9����!Y�׀��f��OL���Ks�.���K�gkk{6N^�$��F�LFAH��TX�;_��hә}@`9�\�{q�w���۷$p�O�� ������aq�(����L`�v,��ï�r2<�~PI3֖a�5FF򢑑y�+�,���������.��٢C�p�b���fރB������2.�$��b!�?��p:%v�������3�٪��4S���m�s�|{zffDxx�++ڭ�q_� &Y�_8�\�ɯp��C�rdg!�UK�����x���$��YA�{["�T�;묅�gP\��hO�͐�ο>D�̨�x�������#�F�A��r�����C�ܺs�����om~�9�(��7����UF�d�,,�������X/��I��er�i�^撖�ϳA{��^,��ȓN��G_�>���� �>�-:6|���1�c������T��Ǉێ���5�a�o��j�/��,��՛�Y����,���~s>k�0;9A�i������\�N��'�C�5�����7�Ŕ�w��@���B�����ïB^E 1��a�Tx|\V��B'�h��+�B�y[�<n@�u�╽b7���
��������**:z`�H82����<	x.��~��4�
��
y� �!���� ��@%ᢟcJR�����\��y�I�Z�c��Ϫ`y��&�/�����INP��j�p�ԇ=�f�HnZe9ޑ�cjʣ@��@6����A���m������v1�;K �^\R���qѵ�+�[��QRR2v�o,��#���G2��ⱷ!�>�^��D(i4q��p�-MKMOߢ���ܟ���F�M���ˏ�z�|�Un�2�jkkCk$��ֺ #�^yY7_��	���E�y�eY��y��5W~�l��
V{ش\v�%�G	���S�1�m��)FT����>�B8��u�aG��름��-��64�'������ub���;ҜBe+W�O�ξJKė�~�n�*�Z���{|����d�1�c[��
B���A���}�q�.H&?�D ����U�	�}�;aR�zK=D�}F2
��09:��L��J��9ޗ����&a�&�V>��� PF��*
��*hVV��t�r%�û��������+tDuQ���Bg�E�3Qs��]�AcN\]�Ή[� �u>�u�d�hV�X��$��E��R�k�*O���3�Vg�%	����o�B&��糯��:�E�4��Ԋ%�&�KW�e�D+\��$�l��%�\�Jz����xO�$���+p���n?7�k��t�8a2w!��F���� ��x����x7Ⱥ᱇������x�zj�GZ>~���+<����/��������*���k���u�D�>IS���0{o�X��p�x�|0]��#lemMB�x���_�\����˷�ܝ��/
BZZZ�hZ���Py̹���7^�_�{Q���t�/uu�Յ�QPSn]�X�Q8���?9�.(�r�PQ�����$7���vB��UĄ��m"9az���E	�cn�=��.���(�b�(p� SaAn�\�f����G\����
]����BF@	��l!!��?�B��[T��>BD����re�J���`�
x>�Ù��|�"���x:��heP�nl/L	�h����4������F�Uuh��,����&xQK+�`�U\n�]U�7(�TN{yy�>6���q~�ʝ�
��!�v`#�:�Iڛ�^�������9)���� �B�����@�?��6�^����&s�+Z�s�����) ^�;>�%����͔�o�HH��9F{A�
��բ��#-R09��Դ��_3Ta��Nm�A	��H@�vp�fJ�DT��M��w���l0r*"�:�XOXǏ����e%�d����1	��Ϥo���)��w+��=�;����#�)�{�+�rvv~�����CP~yh�ҧҟLԲ)��^�
*@��?ޡ�9C+���-P�pҌCL��7�aP�T%s�-z,�^.$ӛ����tWA��\��%7߲G�Ӆ䢩����&-�]��'����&y��`w�~���w8� 0ߢ��V`C��Ph%���;P[o>�n����J���v*��A�r�4�uuw�p�}�r�������H_�Q��A�	Jc豜�ł� �\��/N�w�L
����;t���]1��s|wOP�u��;�����{%����g��rȰ���x�ꕙ�-��;���L�JT婛���ysJ��̱���E�"�_cV��6�;��L�2C9�KEQb�(��%�o��K$0��gx���@�p�UrN:�h��a�

$C���z���c����E�(Bo���g��Fg5=�'�S�+Vz&���t�Ş�#LtK�\$� s{����EYPr�pM�"$�L]�`�)7��ԉ�O��~[�Y)W5�.NKz�)���4<�G��5���%��o�)1�Ǯ�{���pmQeYj� b?�_�Б^�9�_xV��G�Ef����$�0�&�r+�sT�,t��{��b0�s��� C��k�b��b��$��Ⱦ���x�IСb�?$H(��	�OX���P[�<�T�6�t �l�{���;�� 2|�&[AI����k��nuu�끂�5�'k{��o ��x�(�e��0Q�-�z���e23M^��#}�֒����;QhW��d�ք�e҈#u�4p���f��8����5
���G��rY�_�i6oN�x�Y��^��8����)O��J�|��2�����K�@����I�v��=k�º����&|N9���j����B�DI�xB�����v~�8�)��UL�5k��	��rP mO��ا����}nXG�$�i�̋�_	�)�4��mC@��v�a5~e�D�c҂Z"�;hW2�O[��F�%<Y!]2��{�bdj���|�8H�����/K�� 2��}%5��^��܇���ǧ?1%�"����ҖD�m����jؓp��_��W��cB�c�j8y�)�ԯg���4ݺ�-��O�P��L+ΑtN���o�1!������rҁj�͏�
Y2|s^oZ�­�$1��z�����ϴ�')z����.�x�}���{
�B�
���x�PKKKI��K���P���x����"��/�7�N�e�����ͻ�5X�4o���b�����o����Ö_��<￑)&�*���@����l�޼yc\nr��w:�.��'���ND�4�%�A�B6f�O��H�6
��"��rP9��V�4�-r>|1w8� ���4�h{%����1�F�_��Z�QN!��S ߶�U�4Ř� pq����?7hy��O���G�l�I�'Ɖ������o2q�{q
��2?���*.�K�t�Yg�5�U�#
��uI-�KH�q�9���)�T8��9!1�/��,�f��|tP#���vl����/��O��s���(����;�t�w�ȗ��z˼T VH�S�2�{�+/D?݀ka��&N�����%2�1�̆:����y�d�0��p���,�%���L%'��-+_���@��Ԗmo.���Y����ǹ���L%�N\\Roi90봪�*�*�V�嘁1�W�,$L�)��ҒL'�x�i8%�k%�>�RjEs�r�0#�C܊��č�+�g̅
S�:�gx�Nx?��<�vJ��EAs�*����[\H"��9�Fԩ�2L��u��FRX�k��G�+N���D�����>|W���_���-ϓ^!��*�^Ysۘg�N�nJO�	���}�p�z�3���G��C���D�[���ZeI.�|k����@�ΑOa��U�'R�될`׺���l$�\A�����"�� ��o1	�A�0*�0(ݾ�8a���o�7�Y_�8���eF>}Z��;Y�C���aܜ�q/5c�;զ��q!!!9�@���J�'���Su�
n����b6S�Qc�^�}�$<�*���G��a>�Z�Ҕ��Xi=��WW�Ӽ<�:$�<	����!��j9ݹso<�I�ڊ��
7��� |U�8�̰,J�aPnQX���8�aV%N�M��{_~h&\~�F̦���<+Pn�g��ɷ�rj����͹ /�ii��= C�v_�����u��a��ZO�W�y�F{al`���m����*���x�A�С{�F㯫��d_�b6Ҕ�9��������3�S�Q2nx2{�^]�m/���~x]"���ZLJ\'���W&�rsż<b�:��oB�=j`u�&f=w���~��3ښ�FEEթ�m�Kno^		�.h�4U(��$�Q��C�ەg�0��\H@%�Խ���$���h|u����^��z��9�yZ	��^�h:�N�L�����S{��ޣ�+��UM���9���3���s�w�����0�Q�Q=vX)����� j�Y��%oS<�(�QǸ%� EzVT�\����Řᒵ��5yMH�ی�c.F,u4�v��qނDX��eX���|a�ׯxEՙ\��>���sI������,�~�5M?�r
��Jv$Hmy�"^�����sМY?><�q��e>�[�6aS��e���t�r�L/,� �*���}��S;�\"�P�.gl64�ѐN����W�洬a��`F9�Z���.��6"�I�>�i1~�@s���P~�腹_����H�D���ST�r���<'�����Ĥ����oS��2ͷ� �}t��2� )�����o�
��,�𳰱Y��
��G���~�L*�]��}��z���8�zT%���<a�d��{���}������]W_z]<�iT`����(�[���=/�LXI�� |�M�������v��f���x����x�<�RRO�d��])�������K���$qX�T08�\uT\�)j�{��':��ޜp�����ݪ6����r��`�9���W���R��ixh]:U\� �Ɉk
�G�l͙�p:�]y�-�¿�Ilh�}����~���;Kk�� �ޏo����*��9��Qv���^�j���im�O �4�X���9I`�L~u���}�&ޅ�}#q~~v�X�	3�TΑ�@�ͪC�N��W%kD�^�
�m�Ւ{��<ٞi�����㿧V����&�BF�E^���7�Zl��mC.�\�&(_w�n˩��F�)��|�v��[~5�c�l.b���{�d�]ʑ��iu(54��Ӫ+ג���]���f
G1���'X�bd$"���:b����綄�(���of��w��R轜s�>�L��3,�|���
k^�ү�, ��Ə�ͽ�bf���U�It�q����Eo;Z�&�"�&,�y9���6S��}�=��V�|#Rd��M�0�<S���x��F IL����y������:+�<�2G��w�`!'�(��~we��'Au�5���$u���?#�YG/vLG�ۤ͞ˈr��^��dd/!)?ږ���,��.�1�/{r{�]�����R�t-_�Uz.i1M鑿~�SP����wz����+��l�\��F~�Y��s*j�AqI��SGGǵ�Z����7&����	�n�u��c(f\U�El��2_I�xU�GU�:��7�������L�o��x�.��xP�b确|�h��<R��ƨ�(((H��j�[GSI.���+U��Ls}��[]��z���z��\}�ե����ysX~�L��S"c�ӥ��&e��~��6!=����i1��)�1G��bLm ��g��X��'��v'M墲��ڡ����[��| ����D��F�E�WCL�p��7'��t����Pc�� 7������<��ʕ��0�*�����3�9]�Ш�|H
㱼9ٻ��������Z3]��@�Q=�jrM�(T�G�g������,4v*s��+/�1�ox�w��]� �SU���(����g�8��1�D��c�]��,꣞�kDC �(㲺��_A� s�v�@�-���	Ù
bO����a�-���g�r�~~��Ŕ�۾b�u���7 S��G�5���O�i�����^W��~}�+))�L�"K�����Q�mRWk�
�b����p{�6)��Z;FA��e�6:r�o�ǯ�6����5��x�Qg��g�(�{`�:%3֖��"nӱQ��V��oKT}�j����w�
��qdV�.���lZ�ӧ�������2�T�rU_��F�6o����[r��\�}w��r|�h��{�Ō ��tt���}�k�H�YTe'��F������V�H���$��<�pZ�3,�������~��-&:f4�Т�����r{��Z��h %z ��m�?���xy�f���{¾l����;��D!���̗��ڝ/7+Z��BG��I������l�d�!p���y�O����6��Aq�f�^2�l����L�0�X��(���?�g�ʣ _��r�>�O�9�Z.�UG���ՙ/h�ˬ�_���AJ~��JHOMi�D��0r���N���y�BG9s�S{�����ؐ�o2"ݯ7�B��" ���q&��������Z�_����
l�%0V� ����+�"dgΠړ��yU0���D����%��T:�����뽝+������Z������[8��wy�`�TO�M��d5�0~����~��"T�FF�Z�jAk�	�"1�4���q91V���)�e��/�;ȟX���፯���zZ���"N����|�C�`?R�UQ���G��^|N��/]�Q��o��seH��Rߨ�������.4V/��]+���+++#ɃIţUD�^:S'�ʠD�����s,��q���2K�?�����aT�O>��!=�S�H���*6ӯ�	�%)D��b4W����@a�GӀ���P�_�-��R�x{-��߬Fm9��fT���=�����r�q<t�1�Z�W�(�cb57���e��#}�<�ت3��ϡ!�=��c�=���D*V�d�v2I�/t�tm\MϬN�4a/��-��A'������]��8��`q��~����
�����U�sܪ�t)���BO #$p5�!r�GF�P#��P*>?}S��ku:��Fd����@�V0?�^́��N���Y��G;�a�.+�|�,�b�>�t�b"p$��>��թl�u�w"���}�3�9Y�aTrk��v�s��z;����������,Ly��	s�~"��"	�`g��[��R�[�=u�2�e���jA�>;��B�}DX<��%�#!���8A�v�%�`umif�STZ�����JO�q��2��L�e���[f�}�9��f2���J;�R�h�(9osӠ%�P�Ԛ����RVS1�#.L��]c��*>��~��ܰ��xNB|<�潭�!
~⋐�ݜ��� @j������3�5c�v�ݍ��}�s�
(��/DS�:Y:����Jp�RW$����K6���7G�7�,^�4 ����#���N���R��Ӣ�� c7���|��.�H������ Z��E��~b�P.�+88xS[�<�b�R@Y��1��a�>����"�FFc�X)�LS˂&je�B!K&X�j`0�4��y�Z���Vn��
�{��O�U1�Z4$X�~Uf���~�����?�����y|�]w���&�0�Ϝ�j��j��fw�b���+���q�����ͷ ��Eh��D��ޭ����=Y2�\����ӌU ����	`�����c�Oo���O@ZdqDˏu�"��.�h�A��>��]��x�<�vk��b��%ͷ2O�����g3q��1L�ͽ0��� ;{��c���2ʕ�go��1)��ʎg�5LXi��*��폲~{�-�h�,*�=��t}*Ha��?�� �j{���=����N����1c�(���1G���Ӡܯ�1N��opHa���{�
�����~�����h����I5�Q#6�G�"�m��{��`���
F��˪�遜�O�k�5����軻���69�|݊|ז1�g_���9r~�[����+*w�J��΋����@P������m�A��ؼӓ+0=�_�}��BÖ&���HRdv�D�r[�+X.2m�|�r�C�����EGXu�$�A	1������W�\�8��� �5��Jv��Il�3���c�#fPgdp����W{��$F�@*���O��bu��`Qr�>C2}�X�\�=�j�ރO��������V>$$��&���n쬑k�*���e-��n{# ""����"R��
��24�و����r��n5<0�(����'��0E��iV;|Ya�<v�F�ԩ�=�qL0�P��x���e+L��Q�]
�#���
�t�4N�0�4鷾ґk��ѣ�q��:B .�s�-�ffc��l���F�R)�|wE	�X���b�%�E���X�'��\_n��9���8�����h��>���l��
5 �.N��q5����1#@��iQ���0]���̃���u��e]������U��}�C�g��8�
����k�6j����QL8hu0��h�պ�V�s��2m��Q�K_L7����a���7̂v�h�F���L��6�޳l:����oT-�?�[v�$��OC��Q�E�ݭ����	W�ΐ��y��
�(pC��}����`I�����0N��� �|��X�c�9�U
���a��� :=�[sz�iG'�������ԆqHn���~�C��0���:y���Rg��@��{*�O�-b�b����2�o�8t��9��d]0zvq+fzv�3���Wf������Ε�y � ��G|0H��j1]�O�7]G�F��[p٪Kn=O��0y'.\�p6V�����Pb7��� �SMW��F�:�v:�����~M_�0:��� Q��[�m�==�	����4��� .���~eZỉ�-�#�sq>�?wePi��dY��-��*���1q��):r��D����~�2���&J��� ���H�K8�e'V���EE��$=��KT
� �&�M�Cj����`�rĪ�,V.�̷ޡ$��6�ŲaL/��N������uKL]��I�.��'2u�j��T�5��x� �PR]��锇0�G��m��I8��5$B�(����t��B��=3�������J>ʩ"�:D�/Ho�z����`C�̤�SH���2���� Y�|`���㯫1u7�w�?&��~��]m���_^w�!��5_��bdl�	VRk a6ֹs��PPQ���r_ �_�KC��0q�Pk���N �{jJ���l�]�Zz�]�X�O���6�t}�ݱ�f�r���MʑzI:��A�w��vVk0�%f�0o���y��9��
�Q��
�`�};m��`�����Nz�_i��dX`��o�H�+�U]@�SY&}����b��m+Eۅ��&}D�
�7)��!�Ĩ��V��5䲯@!6� �e��Q��W�����Ts0j	����;o�h�¤/���0g�:�0�f�օ�!@�^B���s/���u:�jt9��0���FV^����͆�����&�9 ��I����ܹ������
�ƞ$��g�/�%�V�g1(è�ZC��y��ł*<ٔ*�f�.'��d�`���P=�p�܍�p܏U����{̨/�����-����<�����Yf����N��	���,v�V�j`�.��b��"�m������q�}�bU��ȯ�|��T��(�2
�L�!!!	π��hR݋:�Q��t��ϡ���|���#W���C�-v�`�I�v0?�V�0)u��q
Л� ]�|A�����y�&}/W�Q�@�m�K��.�@ۛ��m�_�{j!Tzvtrd>��M��%�??Ə|�	�za5���ğ̎L�Р�.G]M����p ��_�UH�٠b�4�:j���h��m��d'Q� [1O\ M�y��>E�'��+�/Qt��Q�ިU�"�:�����g��m�xq�PIL^H%W���;ИU�*W��>Z�y�'$�k���E[>�8���P)%����t��##n�h��T�0v�W�iT ��ޡ���B����������_Ek@�lþ|��{�&���ŷ���x��㯶L�1Hw�%�W�#�Ux�Q*k|�����̀���D��X�P�v��łv���O)����*�x�;�1�r�ȥ��>~���i*mx:kw��ڼ�h��
��R�LQЗ�*�I\5�nRN��P!�ر�e�f�9���.�P�������Z�QG��jyN�a�.�)J�;�IV�	e�MI��J.�׹s�#@�P
)���[��}��'��/�Ũ�A��q�T,�۷�Uݤy�\I�k���p�^�����ĵ�we����&���u�T�!�l7�n����1�iw5����pwk���G�J	��e���Q�1�I�!���#�d5Y��xGu��;�a��_*��*t2M�RG��8c�ܽ�2
6H�p{�)F<�$��s�3����q {5H��Hߤ%jE�G �%��?X�o$R<�ؼ�=�=��vg��>�;��G���?+�3 6l�3f$z��cu0@�e�����{�_� �暵"�}�Q+�C���Sb	���O�t�����+'�g���m�>���i֐�*sk�����Y� ���X�3���Q�7<f��Pj��j`7)~��vuՀR���HM@�&Z6��U�����d�=4*Պ�r�kN,�,1�ڡ�gg�};O�T]��y��E����h���\���e;�YUe�\<��rup9w���mRj �X�ȄwV��y��X��)�nW�4Φ�/]���Y��&n�F9�O��S��a��슏�md?����H�x�ZQ�mÈ�����"IQ7���2(R.�Lso�`ǖ��r*�;N��p>�Ú]3�@3���eE��]�f�j\��6�a��(i�V���~xB��J�dߎpcXj3`���]�bm����ΰ������al�h4V�ND4N8J7_,���h%���+�镭J��������Z�4���d{����*ڞ�9���Z�z�5�9��'e�[t7B�o$sP�i4�[�z�"{K+�7�l�T镃�0��4I�	ms��"�X~�?�-'�2W�\2zo\.ր����|p3�|��Y��+�|~��}�k �H������C�z�K�JW��+|���َ}I�:]3 �z{�Y ��������=X�>��9�TA��ʙ̛cT��Q�/;ASc]�5����*���d_�����4��]�Z ٠��_��`���M��������)�%�3��͚�:�Q�J��N���	��<p��&5�.��'���Pe�.n*�o2Y��2�J��������a'�h{�Q�x�xgNN�g�X��%P{�Z8�'�0���;�@���l�:'�~�G�q>׫�}��ve=����|ޢ��r��<a��,=F4%���?�O��������5�q�I�hn��[�̀���5��Ҕ��73����Z��[1r���b���w��R��H�q����ƀᐴE�B؏� ä.T�\��dg?��R�b5��}�slJW?��ym$�̫CqS�7��+#�c��r�c��3�������AVv5�\��8T�
:�"1J
�����n6s�%�h�5�6G��2��`�c+���Wu�^&ԗ\�L.hb5ބ��!N���Ħ�,��mh�ޗHF�G5�Q�m \F8UvD*��#�"Gq𹸵R\^�M����E�)ّ�A����[bą�O����T��R�؃0�� ��~e�n�~ �Ԥ�$=>�7Jܚ]���s��G�T6�}�*ڠ����"�Sn��zh�6�)Q�tJti3��Y��t���u/��\IAŽm�����ޠ��ͦpsp��[QyP��� �(��{������DF��h���k�4�Q�2*v��FI����)�����D�@(>��$\E[�lTD����?�DdbN���)E���V���e��e^n7	@�\�惩��_�,T�wʣ����c�c��O�W���
璹�u��^��(�^�_5H��Bv��&oh��)�+_�������h� �`O��Yf���� ��}.'�܆"~W���C�¦����T4���Ҩ�!�-�,|ۊ�X�n���5��E?mݤ��kv6@�߳��X9>�	��K&O�d��S-� A��o������~)�3�m��O�I���V  V��r<���{hs���G��߳Y�J4�IBB>�
��*�=��qzm�O��q�p�v���a:1��Ou��B�#���ʾ�y�Zq����n��ě~~~��,g��,��-�[2�5��S�Q�V�yMu�ߪy_�}%��__?��$~��3�O�����ɄS��s4��6ϭ�����#I���q�򦾾�/\�,E���G�o|�	1�B�W���~4F�2oH����}5��#x��,Љ�.��(Q�[�T����2���m��\���,��͌�xVa�= 5wțB(�����%MYħ�
����ҷ�K��PTl�]���eA)'7Wl�F)�!�X�챙��[ء=<�GP�D���r��˔ۛ���r�n����@k����iʢ�����}�o/�Ow�GTQ��Tl=���p5�n�w���	�I�ç��J�O7 ���*��-�����s-��ےkc�:s,Xm�^����ݡ>i���ೲ�vmc��+��Zt��X�А?��W��U��"s���ʡ.}��lf��A��E�;_�b'����.R�%+��w��-�H%���<��ܭ���g��,�".�bh�㳒��p)u��n],�vρ��Z��<ܼZ�1���$�5��
�BF����%�|��]_mX�@M��D��o.a�݃�h� ����ҙ:�k�������=#o��O������o�NeE	2B���T'X׀��JԾ[��r�׿�E��V�W۶i�P\UD��Z�j��v=���Ѵ�l���#R`.vj�)˦�q��M^��I�f P=�%iύ2/7Y[�w���}u�W�t�����l���gx����@��8�3�`AJm�hÃ���Ѧ-��#Ӵb32?����� w����wi�g�{�jܮh�o�����E�2=��?�~��I��g�������v	Q\���3e��6�m& j�_g���u�I��\醏�%_����L���Z������6�V�Yr�>)��T�v%��k�P9K���r�3.���l�]AO���ȕ�On<0�z�`�+��/WN��	�}cŁ_��;H\�\�NKO�Ix����N��|�i�ճ�3&F	�p >+K�wm�TEWWw�5J28z�:�	lr�uwX@�g�N�P�B�`�ե���>ۉj�z��T����%����	��k�VU��\v�<�O��F��m�8�cz�g�<6V鐃���#G��E�j+U8�����/���~�?┵����}�zz��_�.��?�:q��5b�c+��;@m�絛��#�r�n�5��:� �E�B�v�������3�?9�BD�	�	&���;}b��P�`���+(+��,J���M���H�tu�"K�x^ɥfZl�o��*>�n.��*:�O+�<��F}�X����&���ռ4�S[��P� ��6LO�����;uǕϏ�g�0p�+,}��4Au����ƿ��1:��Ц^���D��<)���:�����.��'�-kkk}�>n��Ea ʨ!�N:�������M�� ����*�j���2���[���4��.���R�q4fmo.� &޹����u���z�k�F�uT���ҁ�}�?�lo�V\��^&M|h��@d�j҉�=ҭ�Z
1=�_=��M��1����	yK�xYY fh�47��݆�ڽ�3��v���@�%k�.'���o8�7Jۢ�+6�{�wX*ᳯ}�5{K���X37��ڤ��qF2duȏh�:VA�FK��f�3�a�!t�QG��rc���������F� 8�P��l�đ���Mf%��Z7�_�bI#�����z��n�x�3����7���kx��b�u?�Ax�_�!
��0�?k
8"{��oQiu&���Ǜ�/1U�j�_+vǷp�cF�H�8ą|.v�n�/0�n�f�� ��W9:s紹�9�%�S�b#)��%��SB! ��V�<t]is?��]����ǝ��a�wS������&)�V`��b������0O�M?��<����� �m�n��)��>…ח�m"�wu�����=�@կ��75)D��i��@�L~���&�'uF���Qty�mdġ��\�l&gd����/�/Z����@��iqz mA��O�W���os�l�tk��~tW�%;�胈Ҥ��{g�JX�{�����ߜj9�x���5kI�A��IY[�)��%U��h�fq�%�ɰ{d\ޡ-���+Kܸ���*]�T@� ����¬���%lP����8��sߍ��Cyֆ^�I����mp4�4`��r0��y)�	�����u\(�w��YVѹt��{rv��HY3���M"{�6M���b6)r�۲�z{_&zzz������a��LDp���ﶣ�-�YR$}���Py�Da%�����z���R������c���B�/O�|)w,6)�B&F�_7�h������yx'��+�i:I�J���ZP?f@u�ZFO�@	��p7S�}F䵈��G6��f��^TQy����*��*CL#'�KF`�7�P�rd���h�sssO=��(Q\\����a������Je�bs�٢!6l�:%:� �)�[��0�3b����Ku��ak��\'�>�ƈ��wvj�sZ=S�Չ�a0�ho�!��K�,	�픪�"������
_���[��]LMy��� �e���ϖN�}�ٔA��^�4�[�8G�ܷ���_VWW��$�␴3�"G��F����+n��i�3��P��톅H�ܹR���Ӽ�韏�N��%/?��1�]`�B��o���rt�kզQzǶr�{K]a�6���!�{�W��?�����e�ݧ.�r\��� ��}Jw(�3���a��4����t��) �?�T
B�I�*�u�n[6	k��r�?�~/&.N�]�#͂� @Pa��K.���۾�_���F:w1�� ꝸ�����9u쿷ǩkX�3S�y�Lz!����Pb����:�d��B�u&�޲�#G0���W�n�|ז���a�@��a��j	U�-hr��D�y,6w������~�]ܿ����--��z
��֏s���?���:amm-;�����H�ԏYº��~��L�˗�JL�j����Y1:7���G��<��=��6�X��L?#���{�c��V -�Ƿ���mtWm
�����
�|�|��&{�L���soVk�"(��hP����m(D[����;�sp���^�6]u\�~{��xRFy��?s4��ӌ�S��7~�h/��j�F'ߠtK%�i��s�*�?�#�X+��
?�_̾��)�z8����C,�,�|�:������P|�����9��lt�l�OH�����U�j��7t�!v�q������ހ��c�߾y
�����~N0��_�b8�k��}G������9��eq���Ϥ�*��.i"� B��DC�����2o� �?����,^�mb���΍L!f�}e���'�(����665�V��S�(�v� x_ !��A�3�0o!����(�r��x��cP�R�J��#��q ���j"l5�tQ�̲��|�㭡� ��)���mx�k#��"SSS����
5�k����4���Ad|'��2�a���x�gt�ҿ�����}��NXA��ʰ�z��}�r(b=��bظ)CM8W:Xf�jqc��Mq9`�u�Ύ�7��{�
��IPm�G�3+!���WF��4S�R±�S�7;pf�|�����@T�]�!t������� 
��|*�) B�7����eF�&"��D�m��������#����9Phg�Gqi�U�7�E����_N��>��b��01\��<W�g�uf�AǤ?:��$Q�:����ڊN�R$�N}�5��q���Cܶ�ӳC"?������ȥ���x�ùd�^R�h�䶙X]j��}'�~vW����1M�
��
�_��VI�O�a�8YO5��T����^�t�G�����,��?��ß�S�^u��xtpg|YRR �ݖs(� �����^��_�%��2�� �\�i��Yθ�r�q�L5.�?��;�������Nt'ҸEF!��2Q)#m)+d��nJ�*�2*�!{���2:d�PFV������������_����^��5��������'��=���]M�NT7mo� 3	l��873�m�S���"ɶQl�)³���+
c��Gz����n��������|8Q_�'���5���ה��˜�mQn�/
Dfo����x�sUL#/�q9\ktV��~�~%l�s[O�k$�{t�u�g�B�a=��[m�3�*/w@���V~�D�!2Ƃ���5?orq���S����.]��ZU|Ͳ�]���Ǻ� �kl��<�jbbˢ��^2n\�������哌�< A��IڶdڛxN�dZɬ
Xb�r���ﻔلz��5h !�2Nb"X�Jx�
(�����?���a�#���ׇB�wj�H��q�md���"����$�tҼ(�:���?��WP�8-#፠�foewo$���d�C��e�[��3���n�L�������nq��TUWòW��Q�����i���h��pw����i9*''WǱ́�[Y���m`��iViC��'�����
��@�J�,��)@r:B��.zٜ�W��[��L���� -�"�k��5 �������f��#ȔP����X���A:���a߲SbE`ڰ�L3�@p���
ue��XB]qh���/o�?��މ3sΛ�ID����o�#5f��][��N՗/�yQ�}�;�1F��=NOb�Þ��/����톻���w�$��E,}�EU\Y��� ~Y[��?�i a϶<�ߺ�#����A�������������C�1C�yq��e5b�X�߷]��!��L$e�I����xH@����/���wKc+�Gz���ov���ds��G�����w^��G��pj"?ܥS�)����؆����{����roe�7`iy.E�cm9 <J�RA����x땅/�Y�z�Eo�˫�A���ɇOhmG�,�����7���ְ��*�i��ɣ�		!|�}14[�2�A7���A��y��G.���؎�HXE�Z��\���἗��?�߂횔��|��OfW��"�8��̗$�j�^�#��-��鏞>]#��T�7�߱��n��Xɥ~gg���T�����E}���d�+�e)�� b$A�����A�"9|x���6Qp'��[�Y�ib"���V~�m�D9�m�8t����q�t_D������<?�y����i٥@l���x�?�<�p���"&���,F��7����裎ZGöq�J65c��25OI��+���oy���{���b6LᑐY �a �9�������[����Y���8�@"y��8�V^BG��9*��}(qk�B��sK�P.��-f�ï��<��HH.��U!��mZ�~/��[��c,��d�u�`��Dl.A��!a��6b�f�'7�s݊`��%� `-��;��m�ps������4}-@��_���I�C��f������J\�-��X�3lfu�%�}�mM�4��O��9�7>���̀������f �^XR�Ԓ��Ǒ5[�~�$a�A��5+q���� G�~��h_�����ir�9`�Ͱ�n�-�(��6.W��hw9s�+��*H�GvI��u��1��K�f�	�X9G�@����S`p`E�"� vo���)EXʃ@��2e`���� ��K+�4z%dn�M���@��"n�0��ݰ�8�I�9�"u������� �.�Q�.���V�=o�M�����G]�P����/��_1&�?��G��`�NV�����z��`Zn��q��`�۰Q��;��;�  ]�{#�okg��tV� Gks���������6X$�J������tֲě.r$�.�i�$������m���hv���q�&''-{�A�X2�i��zI���/(p��3j�0�,P��`X�u�m�n�T�;@�����vw�E��]�u���7:�i9` .D&g;�Q�eq���RE�7J>Â�U������U��B[�#� v�m�i.ù�<&�������gP��E|eP�ٜx~$�7��F���޺-1+��s��y&��f*$�>�4[޷�IŌ��?	q,E���²��w��V��������ŘĽ;2�hme�S���.A+��� d�p^F�?�n�9N}��4����6! �Y��W\ϙBl�{!��! ��`�
�����ȝ��F� ���En/�*V�3-ă
b4zd,�����OarR1�q�)��r{��m���V��C�=����>	(�9��/vaK��tAW��6�e;�kV���I/�፵U��jc��,�W����z���έ�]1fŗ���)�r��o�����뮲]gw+�{�$.�y�(����@�BďX;/� ��-��P��������"vS#�mNbb�X2�Ī��GJ;�R���(O�oe�W�\��R��	�EH
������+�#~��fs�)}b�pB�M��]�Ĵ��<W�x��&���-��|n����6��}���N�0G�`�f���ט��h�`XQ��,o��Ǯ��8 �q���	+�m=��reHt�E�����Ǘ��e ˠ�SKR�Y�zt�A� �gx\�:����QU��+��
����rf߭�.��_G��m�Q�0��M������ϳii*`xN0^��*M�g��\��������f����
���Xd���N�P\�l�Նɽ�/Na�:r�aAeCOTZ����r��r���$sJ�o��I���_f�i���~�ד���>��xpf��
b\��q����<�`�}��g��`��(=�_�^ �r�|�X�rL"�� y�y,��o��$y�<�F���u�`��9C�ۇY����q�w��#�ns��[�h�6õ[-%���`x�a��2���YzȖ�h��$���K�Pf���d��nZ�ma�2'��g�t�V��[��hU������y  R���پ5n����.Z��ƵM4y��`}�g1-�9s�ʳm�1n��[.���F7�j���0�Եb��"��K�(����?۽ֺ��k��s\0߁ M��+�p�g����q�9i"Ă���\�/E��e�������M��O'%������q����k�u�F�`�F�(��Dl�<"�p] =�x���J ����V�r�E�
/������"{�hlR��c����ï�U�s�{�R�Z����mY�r;Hގ��t�Q����p�?Ĩ�f�\`��g`����R����v�YBR?���b�BtI�T�{���₭��.gɭ9��n<M��d�Z�
���г���lʒ��`�Tkajj�9�d�]�ީ'��RŬJr2ׂn.oX=��������;&\ѿx2�eb�h�1��UR����Y������ʝ��=��[S���c������U_ꀡa�׊ͧ5�{�u�'� �
�SI=�Q۠O²
�+N���(w�x��C���3����\�gϏju=����>�U%���y�޼�s�SG�|~��!wx(���!������A5�3�[�͠�`���D-f=��3���p�*)6A7Zu��0S�B���v�� ���[d/$���򌶞��H�`�Kf�vg�vJ��9Ri�{r�����ui�ery�}��3����'��]*��AF��շ�)0mݯ�$#�+���rV��n�����p��d�o�7��� $U�hdl���T�Q�'����iH ���A ��S�d/��s��=����v����b�a�z��fx
r;�$q��A��$c�w���b�@�� >h�f��������Se\�)�%�j]�'Ԇ�`��~��m�2�p\���&f��փq�0�:��@�X�����QF�4����<��<%w �ih����:��_K��h/w�?�ܲ� fO�����}�-^�j�I�mjJ>���r�]��������(da7�I��v<�w��xb'ytv����V�����"	���zf���Vot��0R�`�}�}�q$��|�%����4s�E��Oy$�bPv�"/؟_���$�K�]a�Tk�]h�Q4��M�>�|����8�����1��?$m=��4�,�|�r��;������pضf 3D�
.��;}@��9ˁ�	dP�_p�G���qy�%�@��sݜM�L��g!��M$f"<���i�l��k��"���s��(r� 9N�AH܌�2|��s�w@��}�d�����DB����O�`�B���_ ��38ŝ����tm�Jk�o}pWl���o�F��e�%%%1G;�o�'���q�ȳ��mBc�37U��)��,Ix�j1:��"�wǌt��T��3NaQ4��O��ZY%�"]/w#�Y�f������'�3K�Z�co%wT~\w
<)V#c�Y�V�ه�/�� ��_K������Y���AT��%_-��'��7�
,��[X�&����������L{� @��5ث���!���ۡzt�<���컷��mߡ�8#P[�Z������/����B�B�1�i�[�����x���IO+�vb%��7��C�8߷|������Z�p�j@�Yno�o{(�e� |������&H��)+��FC0n`�}ܽ�-���0ƙ1vǍE-^��p�;cC{����a�����|��A�����[��s�	˝J��g=g�q��|o_C��om\���6<c�*(kr��R4˅J���d�����ʽ��B���W�96�`�xOE�a@����I�bK~��$.�y�!�����\guI�����vt*,����V�`xڙ�
 �*���0����	}{Kɮ���q@N\8�9��M��G��ͳGr��/*2�,'"�O�؅�[Y�Rq}�?��fQ�#�3����>�,��Y�,�2�f���#����w�?��Y0F���1��hN�
e��[�smS׼�N)��&���lR�	�F���SÔ&�1��0�zKJJ��O�ԑ�G͆���a������a���v_?)��}IW踈	V�S�o,Q�<�Ņ�d�\�g�#���f�R��M��xV��opZ���c,�n���|H�?��!f�k��'�?;��dq��EZ��H���K2.>Bov�.0/;�Ϟw�v�nu�����uO&(�2�5t�t�%�����ߞ>}3��ϛq���:���`�5��R%zUI�SqK�9h�6�3��m�z��n��xr�9�k�f'[��U�e�QvÖ
��}ăsW4f84�a34�h���������+3�*x�g��X^���"]�+�����2�[�GR�V^�l0�.VG��ܽ��m=xT��$�+�ӽ�)�.��u��7��f�TOz)L>�1��R_<)�\��/����p���q�|��ڵ���B��p�r��$2�&��f���[-��공��(�6�����!<� #�K:���A$1-M���&(Tr���H;۶�7p���6��Q=_%a���^�gQ��F4D�0ï̂Fz붰|H- 9�����q2�e"ɬ�v�e��T����@c�UYX[�#��nX��7��#r�J��5s펫�v�!�o����B��Pŗ�Ѫ"C7���ɧ�l��P��r�Ѵ.H�b+9@	��<��G�]P�����;��r��e��lrG�%.C��;��{1���x���oe�V^K��)�TИ)�`YY[+�hŢ\<c�_�mQRR���')���7{zzh��l���pKA�r�_$Lg�.V�w-v	J�V��}U7����9���0��]��9�g�YHp�ucXE�ӃuX���6�C��h��\��S���Y���� K�z�[%�y�۪8=\��gb��˧3E!c�p���k'�]��{���`�.��,b-/����Y�XM�5�с7���n�K����/��.�|z�ҏ�3?=������6ٚ��KKv�l�,�i�����[��A>>>�X��`�>:ߦ�=��2�؜��Q�x�N��Y�S���
ϣ{C�"oX|��o����hvv���� ��mЦ���a^�0H�}��pv�1�N��[�$�ӑ����qd�;C ]mn�W�c̮��~M��^��s�A�X��7�#=_(Ǥ�bM@om�X��jӒ׫y-���l�}X�gp�X���N:�H�Y�3���
�̀'{k��%G���5S�U�� Uy��|�U�	].�5E�~|��ˊ܃���E:漣���������.���va��Ub �k�@�~}ЧܭH�~�sS���S���(%> �H�عж!ݦ<ʁ&Y>��w���ѳ�	��8����F	��b�{�"U=�0�Z7wZ�5�b;�%,���v�y�ͩ߄p���h|�),�W&qO�/��D)'����"M�Ō}�Jg���n��%�(��,TV��l�P�xuړ@����t}�V��w�<�C��a��F��]�`i{��^G�f�y��3�Xע��];�	�*P�X��m�ҥΓ�������	�2����%�o��t���&�����P�|�� �QhI����0�IRR� D�rX��
(�g��n`^��-�n(q�[׶������C�>��p;�B��_���c,��w]зW�%NAp�"���^jO���`f�C)8�2z/4���F��FWq(G����= 512��������r���՚�(;��dNU?���]���A�ֈ҄�R��*��B,�����tNb�Sآ^��%��-�F�>FU)�1����6~�sR�i^�x8��V�=�t�
�ZV��nG�u}��<��|�!O^_�lJ���ױ��c��y�WO��1�
�6�
�O�����03w]�x������Dd���v^�S�H,�!+D��"����7�z�3R&� #�C�o�{���nC����&l��-jx���(P�&��G�s�LhE(n{=�an��B��\��s�i������8�{�U�s�B�̙o��.����Qc��7Jr���x�)e�ں)�ע������[�X�k �� O ��-y8V�Eْ?'7w�Zn��]��xH#�f,��Q��W^� ��ϟE+Y��s���^��="-+�x �Ĉ'���ڧ[7-Wv�GK
	OKMm����z�����W6H��������Tj~��w�306F؄r{�X���~u��V�I��;���8�����)4޸wG��t#51�O ���ⅿ��rd8��-i?Y�j�N�o�i����MYo3c0���.��O��S�,�,�����C�C�C��1,��Yo��_7����WG!�HX#��D��o�ϝhY�!gp'F���d���>GX���2���8`�y�"�{Sk���'U�5�ɒ�@^�V�f�Hٯ����� %���*0/߰�������#�����h�%A/��noo����D�I6'�C���2��X������[��F�3�+�,# �6�M0��Ӄ���8)���K�
�����Y��n���h��N�i�O1*V>#����=2/-�{Y��7�nK�&v����7_=L`�s+�S�P��L@��%��C�����w��#ccv������jR(�I�iWe��4mś,�?"oa�P֥_�&� �e��瀋;&q��q�t.¤����G����K&'������M瀍Ð����̿�-5I����@z;�B����5V2_��D��0m��Y���u��Yr�I�����#���1���rX�	���-�ubn�~fp�m��H
�w����(�6��Ç���ʼ,b>A��P}���C5V��Vk0ZY꜏
����nD���gZ�d�r�Nn����VX�p��09%�����6c�����*�"R7�3sc����-�N���ܙB?t��8W�d�NdH�w���Q`}0N[!��8I��_|\!A��v|���*a�"^7Z����1:s�3�4��������ͻ�6�W�o=:�9"B�ˉ�"jL�y��0V�@S�tD`�=K��վ���P�cj-m�0Λ�������:bªw,���Ŝ���f:�8��E���`�Y�#��	����H|/��m�%���mCcGP_t������������\o�KPͥ��5�6~�ؾ`��w�L���w�d �}��E���>6X)��v�:��bj���45�Sb�e�źA�C4�O������f�қ�f��=;!{�H1z�'�����~͸�����t֥���[�|9|���[�X�`��� [ ;l�ٿ��;�	����!K7�'φY$TW5=}���?	�Hj���&_�7��?�uy�;��u����,�%|o7��!1��F̓w���Ɩ����j��c
1�],��ĳ���9��̼8�0l?�8����&_v������g�;=9.~'<�@�L����B��kbkiܓ$�KD�6�.|��s>���СCU_�� gv*��Cb�I��-X���E6x@k;q���4��z)�kh�u�f!,M�0[#��y� k-��M�M�#�U}C#M�!���k]��v�2KL����+[��5���[m� v���((�Y����g�nfee�!l���UpFa��(�e���||=Pn�v��	�o�����)z����x������a�L�x�Xl�.XX�'b���:�I�6�j 
��`�SJ�<��"V��+
'��IK�wktM>�����[q�0b'���'����W��SC�5Alp�t�R�Q��ފ�a��r8�@�,�%~߰CW�y�g�Fu�'> Y�ɳ��(�LdM����h]a���`�ӌP��~��dA%�h�dBo;å��:��2>���b�DCB���a�|��щ^w�6?7?�<v��������GNo<�"��1�g�}���)@�!��	�ݱ>7	�h�ӎ�::�S���f��z��
z||<�}������Ĝ�#Yc�j��]��%b��qZ!��6�_��>�o��Y؉��  ���7�i\�𳳤��T �Bb���b2�2f�-Ţn� hoO	�����>b6Bo�>�دZ��� �<�l�5����M�����U���g}�0�K؆� �.�k]&4Z��Xr�맟¶߆`�� !a�$�_��^7��"�`��5ӦC��2e�� f��1{_��cٱ�[Y�D�̨�$�;aq;k��]�M�t�M8�z����蝶�oC��U���' n�XՈ�F�SJR��Ʊ޳�����^6С�=�ٗc�DIo"�%����t��.`���s�:3֢&���tgH�B�Y�������O��G�$����`�|����_��؞H����(de)~���t
�WqѨk�-dY(�^v(�Y��ˏ�0�w-,,<w�<I�K��g�m_����, �!v��&tau��P`4����̿M��Z`
�3����{�ɻG
��
	9����:�%i�Ԁ���L�M���"�K���y� 5<���(jJ����y�|��1XN,��x��E��$�û#c0�ebN�B�M��bj��lN��7�+�A߷���X;D�����ـ�7^;�N�G���UĜ;w�E٩�K[K�!S&O�*��Q�t!�i|i1�fؑ)S��6ȼ�=L�`�:I-�깭+�7��W�ضl�}Xd�> ����<���C��-���Ϥ�:�<��M_�S����y����O"����e����P9D~�3�^I����c��U��!�d�k*��v /���to��J���6������G0�s1|�,��ы�[*��8��cb���Jm`q�G&ff*
�LE�_���������������ijjb���]��"z�Y�HaA^60��~��8)�N�<'����z�zm�>��b�"�X�wv6��`�>��>g��<�_�cͲm�ǇZԐ�ު2HҀ��]d���5t+��Q4�/�dg���'���!{�G���α�Φ��v����|��M�68��q���Ǧ=4V�{�������TｱM�X_n�r�CW�sۍulD��E�R	�P������"�lD����7����B���������K�!i���_�
o
�����gZ\�Ȃ��-V�[�89��l<U� ���.�jf�,�1��k?(�@���:�k
X޺UN��W� �N�A:�#��[�XpC������<v��t�f1����OȾ�ƭH��E������ၤa-9X0jǃ%�Z��>׆<A}��D��ra�Ss3�ᗝ�����L���ڻ7�g+�ף�,%,�A�$"�Wlw���q�Nw�2lPۋ�,�驡�d�dG�s^�稨��6���A�`,��
)��A����X�� ���ߪ]W�����B�c�K�3��!2#�������W@�5n�p7w��a�����`�}1W�}�#Q�}i�▘#��� w�u��Y�3Dś&mf�B��`�v�ݕ�{�&�za�bG ��*؟;�%�j#<�#��߶i���/v�1��RQ�E��b_؜�YS�s�XIN +�N����~bjU55��N8���{�����d����c4��13q�}�ƨ�����+���L\���Y�� J�$9������#9o�տy}�����1��$+�5on�eR��̓'��>�ºj�:r(�M��㴓kl�5b/&��������*O�������jY�*	f��U ���Wq/qR��+���-�E���WQU���^������[����R & [���<))����1�ha��b�Ӝ��E�����HKD�f�&
ћ�jz&�X.�7L66�	�)��	�nJS9n���&P	���H�>������iR,��91�[�mk�e�ʰ�+1[��vR�@o���7�Y��L/���?�eI��^Y��6��@�<B�r#%�`_+�����h�(�~��o(�o��&����q�mo_�zLr (�]e�H9> �Y�[�؂�|�n�?�
E+��Q_��j4v�E
�\T�8m��M�������2zLI�#,l}s��7�.2�v��  ��ș�%�2�.*E\)�א�&Ĩ�W�A�jy-|��'~�k�M�C���q]?��@ mk��}�D�n��G�.omu���<�m�����j2�&��m��'�+R��"��c8"���&>~|�)��)K	.j(O�?:^�U�{n.[L���xbelA�B����5P���M��`��m�hÑ���O���k��صP��Z^Ha���Z)���踫��ݒu�?]�c�S�Q�ظ⚨�9l
���F��Jc2b5l��6��������4��Dx�C�k�h��C߁|������gA"_��}�l��U��P�}���9n���?�-Z�9x.%���K���vqV�OWȟO��1{Q$*Lo1١|_�͑��l������Zi��o�����"*<�#h���'�!o"۸<y���L��@���F-�σ���JO���N��D�DM�����0�H���D�L�Tf�+�B�H^n��X&[#���y�!;1x�_Q�Kj引S��Įk�@�������J�վ�Z'��/v��ⷣ�n�*���:ʃ�2o< !b��L5���؜�w����ܕ$-!�h�|S�6��D���̉�R�xi����Go�N2�1]8;��x�-�`�ٜaw��ׯ_o2/���g#|�h���y���O�f��r�����i��B	�@�B���m���M�ɚ��F�e
�#�ts���%�᚛Z��qK��>�(���٩���%��5,�6[=��ir����K��AG�\�d!�?� ʢ˜�l�*���5{�NpQw(ώ���5�;�vj��.A�)��=М�N^s���0z��l�	��85���_�}�� ��u�����4!_�aP/^!ٛ�)yJD��t=I�
�`���T�oɷ��ԧ�#P�hh�p���(��zbЎ�����5�k��G��؝�|t�->?T���Շ�`���;Y4�\�1+��h4�1Z�HĢ�^1��0o�<��5�#ȇx�6�_wY�x�����$c�1ε �yZ~i8l;��W�
���݉Gd捶Ӿ�bљ]�*�����!K�#/Q�w�y���x{A�d؞@�{xp,���޹��A�ͲG_�U���[��Đf�5�����;�jL@..W͗=�������VY�@I~�;�+[gu�4�ώ?�)ܯ�j�5v�[�U� 0��=��*��1��
N���έ�ܬ����g�b^��.�=��+4;�"��?�>|�VS�y�+��-G�\���nb�r[��G�c�@�u%�-	���AA8S#���73�������K�L��I$c��G��8�Lb�S��a[N�\���>b
tش=.ΏB*O"����D����|�����/�R���#38�6�}~�Y����Y�;����{�pp	NN�+W}yZK�*Ta�
0O������ă4=����1��L��(L%a�kn`kX`�@���cf�5��Ɗ����++��1���:� ֮�!\��ևl����=g��T��i�5�9�84�gY�YZaW��1���1�0��5�OX��,Sk��;FOw��z�IՔ��>�xV�i������4�O�cC���U��#=f؅��D���_.��+!�kCn��_yIS 6)��������V@Ү���:K�1�f�$�t>�WZ�̒t\|jI;:!{�x���0g�J���X����6븾X�Wgy�U�䣯ĉ���N�����$������K΀ǀ��G����X�X<�@����}3���6�zMV���h�h���["��
��"k��O?3r���o���?�"ǣ� �2>��/BT,��C~J�����7�*|��V�j�;��m߂p����E��YG?����S�5�1����G8r�	5R��+K�M�$�MPs���&� 1��p��`+��,�&Y۔<{E:,U'bT��M��#6йe�Y(z�לd�$D�pʌ��O��m��]xC�#�7��p9LK��Y�½�Ϋch]�}/N�K(�>�?D2�/���a����z���m^�?13�H%�(x_��#JT,�&�7��k(��|wv�+��ޖ����(�^;�Q|��x���e� ���o@l�vP�K���
"N�#�Q��.�6!��Y�<&�Ϧ��z�'3���	�ds�ëA����j{=c)��N��2��&��>�ii�e ����o��*����{r4_2X��a�LlwL7��cњ�Ųe��22�Cx��8+iS� �p���WĈӖ�( �M ��*M6�w�T �� p�4��H�z�D¸)�#�-���K�(>^��������ױ��ľ�&/)Sg��� �,��ӄ#��=H���@�~���e۝m	S�V~�����c�s3M��-HT�/�0o p�yn�ee��'�qq� P(���5aw�.�CUʴ�5���M��y+�d���X�&8�+c��͔@s�Aq�o$	ny�X�i�q*!a��Sޯ��7�������<W�9[��b���1{�	��aj�V�*Ƒ}�MG�^�j8#�5���m���{_&�7��K庍!׵V�Q�g�h��O-��r�"2�#
~��_z�^�������h"#_#�D�K�z�]o!�5Qp6x��[77�"��\�"�-h8��Sw�����C��p==ZϏ��dKV�!�A�s<�jǰ�O�;�vF�Y���G�!&,��_4f���e��>oiys�G׮�XLK�l���+�V���!ͼG���ÇϖW!��|OB/#���|����ׅT���A !��1~򶁝`I��=�|$Kڵ��z�g�"��+r� �	�řX(�:��J$ xvyxx ����Ft5[.�ɒ{_~$I6	߽a��8h-`%G�6�uF{y"]*	�������sDFdۀ<��^�.�7�a��<�����8l %�6-f{m5VI��a2V(Cxj�����Y7m���=�W�G.��Of�#��n@DC����=����߂ɤmZ����:�8Иu��6_���S����G�f�w�Q승B��ə��˩�����_$����٘�@tJ����Ċ]��K��0�3۷�T�,���}�첝1|I��� �qa��
O�pI�1��b��V�H����:�y+<���u�hU�K���'���ޤ�-ҝ�)4.":H؈��?vl�����^d���}�Y�lQ,��6��m�?³���eN�!2�mS-s�x3�|I�$�Q�;db
���6��eX�K��Ъ
��h�2e���x�"�� ��=p��>�n_�MLā}��o{�NA�q}ծ���jP��8�!		VR>������3M�Ur��&_>F�nH4��cv�G��Z��ZzZ�Y�h�4�(��[ss^R3��GF�������gO�~mꑛ�:\��_ݧ�>��_JByìɱcQ3��Q^Y4�+P�0m5eT���Y�4[��he��T���z�1��qb[�U� �m�8���1��(�X��~�$�Q� j׺%�pU���6��I�-�d��S��/I�M�l�ÿ�ɼ�����V�Y�'<�Z�}'ܕ\G{':�D�oDؾ�_��JF��V���Z��$�����m4����4�ź3�8~�V�X5N�Vh�sP|Ȃ����G��$;���+s�Ư��^�j^�{���ٵs"N�Ui�Cݧ��E_w�~r|f�ao[�<n�(������p/z-C���5k��F���^�$��o�{U��D���`Ll�pֽ�B��z���(X�yD���z"��e��HS�)����ؖ��Jy9U��X�q��	���륯����{���*M�b��K5��\ś�p���n�٘�! �<脒�c�?=���`B�3p��G7�D��ש��5��GV&X���|Vy�>�0����������Mmci7%/�Vf2*�y)�3 ��0�/�b����1��	�V�^}�mA�s�3�+�Z��'�}�W3C���:��Kj���r�շ��H�/��C��W
���N�g���[=�u�j�:4�w�/��ɩ_�t	M�-�Ug�H�2-#������Ng��esjՉ�{��O�G:$�#O-�TV`MN7����Y t
6��p��\����-~���,�.�I�MɋN.0�h��m6�nK}t�ԩSU55ܘ=������f�T��P�,!�W���'�d��HZ͸�����Bg~g��1���"D�E
@V���_&������}������j���丂5��}2��� 0.��pc ��(�����S�H���wq�[�y� ��3Ϗ�G7�Sx���������M/}9D�b��[8�L=#Hz���sY���V��v�`@���*X,b�-�����-n��smZ��j0��Ѯ��S�ar6�}9!20�n��?!�wF�mb�܎��VN�}\l���pﻊ���X���M?5�+��6~���Ma:7����8��b����̙3UUU��c5�p�3RC���-zY���Je�\8�~��ݻw	_p�k,��q�I�z=8�5mqD4��Z#����Q�&	rQ;kr�
d���b��8h��ǃ�^7�����|��hU�����.X�J����|�qN:���cP����l��T�MZ�߉�kj+pdFV�q8F���r�TU�9�3����T?S��t���g�[ϭ���E�!D%� w�om�}�t=`�W�t�n��u�@*�}��PŬ(�)�ɺo`	O��EV���pom���g��+=�:՛�V���Zk�p{�� �%�f#_�Osw-�$�>Э�����E�����!�>P�����fgH���x�$�c���my���d�캺`~���F��Y�~��*K�&�����nMZ�$.�L>�J���<k��h�\�/ �A� �ɚ_݌l�SA���g�@܍��U6�e��XǛ�m������FUx��4������7*c,�����c~�+dO���A�g^���f]v�<w�<���"2;�`-\g�'`���JN:�,��T��,��2<k���ft.:^=M} �	�!�a4�#K,��	G��b�ONr�R[�S��8{���������vR6ǒ�-D�'��� T�k^v���Km�D;yױ@��=XP���'&~lM(���5ãT��/z�;�m��r���Q��a�b-�SLS�p�	R���Y_MW�v��i�i�Rf���@�(̞c�����Tt6q�a��� ����ϫ5� (�� ��J�*Wn�0��B�z���d>�Q�)t[wl ��S���M�CC�,"�.� o2|������OK�X�u>��o)��2���Gk�����\Etx�2�8ҏdڝ�Mp˒t�����:���}>�ȣ�3��1�d=�WRV�D�+�8�k�;�B�r�N�!��)_�ޭ���[{���n�8eW����?�I�ک��n��&2���m��H��,*����j����X�e���83Sc���øv!u���=��D+{�-�Ҿ|ϙ�_�q�p;���v����y�3q��+��po��<�tg	��+����B+\Rb��]*��m%F��ޛ}�>Kp�8�a_ _a���ipn��Y�U�_Y����t^�7��L�B�r�#9[6��#`�Q��RWM��
����]����2��Mǜ�xW���^qı��yS��\\U]}֠�{�� �Ie؁8{�*��7)�d���1>�`��V�8wk��~��<'�(j�ޑ�ǉ�ͣ�[U��4�>3z�>|4�Mï��Ӏ�28��Ի��n�]wt\Vn=��@X�S�S���]�Xd�O~[51' 0��޿(�=2�,�����8�'38bѱ�������&���� ,�	��6�א@�=�_�8��j���з �u\tǮ��x����'��a�	Lcd��7���C]%�hwZ�4�Jl�������U�U':�m:���A��#ёUXX�s�OuU<��/�A�Z�N��'�
������G�b�A%�+�����zl�k����u*B pd+9�a���b0M�h;�"���7-!j���kcE�q�S�\�{r�D���#F��`��مp�3`B_�ّ���7�Ag�a=�2NX���0J�.��n����
�� �L�vrt��s�7!!�L����GO��j�w��*����G��S�H��Zg����7�d��-�W���8ȟQ��?��(�^�h��s�<Ͱ��1���w��tkQP�Z��r�X��3�^�\���}qG�,�AqЛ�u�w{ '���/�|14_XIɪǑ-�2��"���۪a����u�D���(��qx�������g��-��71���9`�|G��	�q'1��*�;j�X��}DE�Y�x�^տ��9���P͵�OGbr�����|i�Yv$���?�E`�Sڙ�4W*J�m��?�]'��!�Gم��P��������W)Nr��a�x/��c��Btf�V$�f�����=���2��o5O�מ'u� J�;��d�G���9���yĄt�G�b�}��[K=�Bj�3�074������2l
���d4���U�X�6� ��c��2M���[�0���V\�K�����uV`�&�����[_�l>��c�M�Rv)\ު�?�5׼<
�m�eѱ�x��MW=>p��u9ފ��	  ���	��"Ś�;���+z_����
����W43t�H���{����<��F�<�9ry��"Б ��}�#|�۷5��e6�L`�U6��rƯ2��Ba��I��\TY��}.��c�!!����k�
��M̀%�S��t�#z����^_��'��xzI�aʱH�>�sltcm����h��f7�ϹX�jY���
@YK%;�Tݱ�D���>Upۖ��l]�ǝq
��|��l�Q�8p�V��	�c�
3ۉ2�a���+�F�ؔ<�w���UI��Q�l��=I�]�i=�~�rhD�m8�}��e�4���R�Y���`��Yc�0�Z�|ѱ�P.�������\���a���`�$N*Iv�+~���O2<"ƕ��	,�(�Gw<�Z!�����[��H�Fݫm� (�v�dףW5�heQ��4Nm�s�Ӏ�S��팬֘��(3�l�Ͻ��?���_O���뢒P�]O!~�D(�iU�lm��O��$kpn)4?'�>]_���>�g@"]�1-)v�Ml�C����M��nQ���i���5���*��}���#A &�q<�c������zk_||�����'�ET*����{�С�˜�/�W�6���5�H�Ư2\��@��f�sѹ��Yec�4�^ޡ��6OB�-��e�$�����Kn�!Qn��ٞ)w�W�꽧��ޟp:�47���XJ������^�Yz?����i�{�fV��YWG�m�1ȷ�ϟjzrh*�ejj6�T8�`�ɺ��`�k4o������׷>�V�\H��VN\�`�{ ��<���������#���s׼Ư�w��Ͷ�	755Qwm���yꑧ�P�)o\���ܔ�܀3�M[��
+hu�8��W��v3K
A/��!�F�x�✍My`}Se�,���Q*}�z6�M�O$��X%R������O'�1���B�g��r��Y������E�����-���)�Zt���̡��"5��¿�UB�Nl�^�p!7��>��gcc�z��#7�/B�P���MX�IAG�Y�k��>WW-�ߤq�2��Ӳ4�]t�{���m=q.)rt�6�6�����!X�<����/� ZW(x�~�
5���"JA�����r�7�-�526�_�J�:g'"��KW��{�� ��[ZV^e؃0�Sm��`�}����o��sĩ��)�������ϱq�h��w��WH�S���*�D�;oTRR�~�E�G
���Gʴ_�ϱa���&ϩ>��Y	Y'�]%�#�D:5��@Y+i8207��,^�_Mq:^�ݗ���5}{nq�׬Zk$@&�SR]�[�ý�`�+���5? �j�nn>���h�9V���+��\��)g{����D�����t�P~�15yq��3q6q*�����ߔ6^��띛4��rhɟI�U�q|�N��E|f�.�G�X�k�;��PǇ�?x	���rg�~���:���>�<H�N=(6��pSWub-Z̜-�6�Ś�`��x��h���.�6<���ZԵ��w�����u�}��q���Lʯj��ͽ���)B�oo+����9�(ۈ�8�YႬq���B3cca�s��_���!$���L�����&Φ��m��XAT���Ia��~[M���"�˷���7��&��T�%�T�؁���V��s��͛ f!o�-��s�s�۞�"����.�'�}ix6�CB�IX5���EE����H�{������C.�c�m<�Ԣ���[�cCv�[��n]�
����h����ا(�U��
��v÷�O,jEڇ�`?��x	��NY"q�ϩ�9Uqqq�{8���Ak�N�C=	���V~��;S�u��*^�������m|�O&�(�{ju���vn�c��a..���9[���{=ǚ�:�u�ނ��ҟѳ�^d�n�g���>�����e9���I7�ʘ���yD�j�&��R���X�ɯF�이��zq����GhM����k��v��� �
�	��Ld9yh�1�C���,$h�x�M�������ȵI����|��c�-%�xӔ�
�r�3( .��Y>o'�CC�	�6<�1`�����{��Yd-���\B[t&�)�4�H�qp�_�؄���M��������G��%/[�!`���$��;!��#�ir4R����G�gk斋���������`S�L��MsĆ��#�䣰M`|�_�^���o�V�:��S�������jm:���3`C����,�ϲS�h��$<��AC�.�Q����������r�փ�x@� ������H�(!H7
��P����
Hw7C�(���5t��{�s��\��3�}{���
�`lf�XXaY�V@��'� �!y���Ut��/}�-���p����K������!��u�z��KV�_���v'�`Z'�n8�]��gbȇ#���'��,GE�+R��a���[o"��VTT;���	.���~�1À���%f�+��@�����
��g�XԄ?��Lk�h�'ݿ!6pP�s�~�D<�m������,--9-Wn۰?���ü���q�3���1����T�a��VX␘�h=���0r�M�3�()-(O!V��m�Q��.�j��a/�G�>���LJg�1���>�W8���+U�b��y�'Vn�i'����!�{�����,�t.�w& ��@!�������Y,�ޟ���-��MBA)mE`#'#�2������T���`���`�5H�p�t!`nH_�ar�/���6��X��cggw���5l�djF�x�-�|�� ��ky��T�)m�Jg綫�]���!<���NZZڜo����#N�&ff�c���G:��̡���H��BP�X;Q���U�N�хr���ԝ�@	G�La��t sFGc�^k����Oi����u��n��M*_z9Uָr�9��ju��sJ7�V�a^}��(� ����+"��bc�b�m-��y��m�NLLt>444�cs� �9L�3�'����4�J깬ze��!>>~g��m�Y��V>�|�GkC�;::¤��O�V�4`�
L��T���7����~��i p�X �HD��W�����֡����3 J��9?��h�ͳ���3HV�B@�vVj�~�#pjǕ�[ew$4�|1���
N�A��k�O���
G��ɸ��3ĈQY�s:@�Z璟����M└�--��y?�wXC��<�ŝ�������ٷL8��];����]���x�-a��l�3`�	8�LW6\��}8��p��R�D~=c��qSS���12n"�{���}:6�������4`�H�m��#����|�R�-|]��@���H%��ċ=:z�f�۰��y���P"B;�P�O��V�N$�~C�G�7&?��#�o��'L�0 R��.��"�dX�%���N�)�H�'��zol/J+�H��TT���9::�+0�'+6�ΩS�x�X�D@�Us�i��>��р�����j�w�a�!<���9��)�0I��:���.�ǲ<���L��������}�P ���aRTQ��VE�/�G>0@�0Jmoo��cutN+8�Q)�6���;5v��D�Gݿ��LT��[ �A�W��կ�pӸ��1+>�-�hZ�t "�?�⫻3�3T�37B����{	��a�,r k�3O������aN�����)
X&0�a$|��;Po�8���8#r�OAfTU�Ʋ�>�?�������fV�oJ�'L�C�h m�~�C![Ii� ��=�zk��K�^ �(�+"D�����F�*��p�p��r�0�j�͏��R �`���L#��߿gR�k�.�u:N1��
����W��Oa��2�n����2ٳ���;��ȿ, ��`���r�z��/��4��KFbPK���&�:�+��%����W��]�E�q�z�1Yy��@%O�Nq���p�������b��vN����lh�������I��(���/�p%)O��r��N��a���L��sd�`�8�y�=��]��5�Y�sK>�9�-J�20Y?ZB"��D�{#�{�,[2��z=�d��� �E_r��oA��Xn6"<���IE�M"�}\VeWw�Tm��8Y���]?�#6ڵԪ�zY�T/���񈄂�Mz�99$�s��ί3U~����u%&f{k�LW����ic�{(�ND�"k_�jD�B@>���� �X �5Pa-+�X�-��,;��l�������D$��r���H*��
�$$$�4
��`avլ?���SBh�"�Q�����|&��ک�t���������Uڤ����a^?�ۍA���-жBfj��mt�i|��9�^�����n��Զ��ྦ��@��mnn�E�yZV^��
������|a�N�Wj�"�& @�.�a�)Z������A����m��ۼԜڿ����uv�e�e�$Y)�P100���1 )�R�����7k��M���8�Nԯ� �C�Tk�la�Y43:\@�(�a��S�%�x,~��t�TU��d�Xä3��:��2��̜C��S���GL��܈):��x����ez��8U���{fvv�ߣ����R[8�I�)	�S� �NJPקR�ޜ����y,��% ��xaGCbr�f!}����>*�JO:U.���+GX�>;;�xEz'��Y�1]��ңE�r�̴�2!d݁=��{t�/"�����P`�m*��k���[���`~��ax�J��(3QwnZzz���Z P6g������*� ] P�oD�->gY�
����'~w:��P�����1��a�Y��Na��s�Lr?�/�z69�_`�3�6��],C�Y�����[|w�l}S�-���O��A��x���lR�.���Bv1�q��L֑/�!�6��vE����6+����5�c��A��H���W��$�9�+%7��7������7	����&������j8!��.���I)�]�1ә�+��Ǌ��ʣP������?�?���&$'Oͯ6N��z��#~�a�As��8T!b�
�s���%����y}F/�e���ש��#uͤp��eeekIEۼs�$թþQ�:$�m�wo��ѭ�L�ڴ���i%�hl�5\�d����"h���@��%Y)6����W�$�\qN����PzH�:�����k�x�3����(���;yD�hi;��zݺ~�:Ͻ{�X���h��6x;�c��1�7�F�|�hOo�^4��|51�z$���=��N����#�������llCT@�ٹ�ڲg��SU}�p�/weN��٢��ԂZҿ�=c`EZn�t6�yS��8i� �������zYج���d~��� �]�/ax�b@���SH?ņ {���%a���xI^V�����:�Y���9	����'5]���C�C"�Y?�C(x���:8@� H��l�L(����e��t$�c0����h��l:̖�ѳ�b�	z���Q��j��*xcaυ;7`ۯ㏚H���*����B?tWP������K�z��{��>��c�����Rbj�-h�ٱ	�J�3s'DD�"�&��?�NC��c���
���L��9(�p\�b~}X�'�<!�˺�8.���5g��療� �3]�vq��/Ċ�lpY=�ݔ�����3X��}l�2��JI�b�+PV^^�H��o��������g���j�O.�5p7��$tw�H�{=)n�����UՋ^k������[��W�[�b���RR��a���(�FaYSSS}�`u.�w�B;o�Eᠽ��>u�O2$e������Z�Jm�a��f~���k1�a�5�b���&?�����c�!<�6�qW��-�סe�W�n�1	;���`��/9t��*Q�ӟQ$���W���yN�3<����1�	�q;�-a��?\EPU8^b������b��PbT���_����O������;,��W�<[_�>G�9����|��uƱ�p�Y�m?x,����T�
�.x���&�=z���gM���F��(G	X���!<�eq�&a,��1�:<� �Ƈ۰�3�4��;�g���ܙ����Y�2��* �P˞[q	0��vWX?��E��]V~�wv^���k��$�z��R�A�C���I�{���
S���u2�\Y�9�i/j�~TS��'U�a���ЈOL�N<��� �wt�Y��
ӊ�1����h/�/�Ǩ�ǏN�Î��%Bm,����+:�3Tp���adؽ�����$nԵ@Z�����ԙ���g�3~�N��	�|_��*��|I�����>Lu:��+%�*,����©n��lW83	�����3o�8��Γ�9�=���X��\g��@~xs������|f���,�;�a�ժ��\���d��G{P�L˙�Hƍ��$ 6z�_���������˷l��7rez����W��`L�"d=$^�s�ǟ� �
8�F��`�޷�h���ׇ����F��7�����ycx�_�Wp�`���S8;��}��V,�຿u��&1��{�Z��y�N�O��)���rj�\ ��xex,6PX-��#a���T��/�J��|W ���C�CY��^L���=�@Y��`��+lX1x���]��Ă3�]a�ΉSô�AŐ�0p���3gNA�a`b�'f��r���p�p�C&8���u���zb!�������1.�N�ַ�����J��7��������_��{ׁ�,6}����[S&��$/���"�M�Xz���D���o9�P�c��������݅���,�
�ӲrS���~�S�vH� \pZk����q���-Y[ �U8���6�5�������+K���w�G~W���߮���N�$T����Yh%��l%�O�5	�0�l\ �>*��� f9~�"`�l(��󾡺oXU�5C�q\�(=�!$�PJL��Țd��q ��R���6�������Ϥ����(U�������B�gL�T����m�	�=l��+j��kp��0���Mܮ�C��q:�Ak� '9����bq3J�Ǹ�k����F�GxLͧ)�����$qpJ8�/.,�g}��m�H�y�B�u����Ny}X�(v8Q��w�=nΩ^�Z �綵��&x��P��lM-\=�HI�z�٭fО !0��7�c'>`���\����0b�#�������6x,��c���XT��mB�FI�:��WZNF@c�oZZڇ}��&�����u}CCe*.���4���ީ���-_*�d���h7*�C^����e��i|�K�N>~��S�����������VWV�>�l�'a\��\=�=���j;���X8�Y9�8�#{#��NY���z\$81)������˕ۺ8T䢗NQy�b%����Q%�~��Emo�l g����؞,+u�=Y
�L�_�<�l��]���ן=�����\6W_=%���������ӌ�:>>�
=-g�B��g���J��v����oіj���9��`������b <�NGZ���QTW�.Wp
�t�YFfB~�(��BbN��LWmT�@�HNf�����rh�J�A~� ��:%�W�!Jz]�?0�veL��9]�h�s�0��3	�c�z�����x���-�a��:P�3�:�`{l��a6��:t��Zo�D�2P� Z�0�FR��!��ԟ����ꩭ(�|.f���74��YWW��=v�t-���mŴۇ�O�VO����0�{z���:
��Ʀ����%d���y3�?'�hvA�w��˓A����n�KK�H�6_�njZa��H�q~�pqN��f��!o[$���nL]�Ğ�wZ�R,�k��s�sa禼��2#����9���~���)y\�v� =�K��n�h�a�vo)IB`Ò6\݁#�hJ���Ǔ��F\8��/�6y��>^&�l��RuSz	�QN=�Sb�[W�r�m������ws`o���VY������R�w�w��ϑ�=�����ؒPst�f���Z��]�h��+|	!���<�Ul���¤O��o�6a �۟�NCtJH���P)��Dڮ�v�vKK��J�`�y��������8%ED�R�>*�cbd�]�Y�}�c;'�î~��z|�4`vq�DJ�Ǐ![�ṺX��5*�3�fE$�N��̙��mhh�\%���T-p}�������O{����C�<�/u���TU�V�UT�����_�D<Z�i'Q�E�>�O�����ߝe�%CXT9�%�����֟��J����� �Ĵ���dkL,J���*q=�(�OK�I���ʟ�f��&����P/di�-�<G.el,%6zqF��~��<�u��`h�EԆ��h�+d��~<1=��)�q�g��6��01Tj{J������k�����fw�z�1��X&�Ȉ7]�fv:�D�iVU���2�.*$U�:� 3��G�D��8�E�,�\q�%��9�>�W��mf�U)C�{1���A�E�X���XH�P�B�S�`�&�]����,7��+�5�2m�"��������I��l{�t�h}ױ3	"|Uű�J;n�e\d^}B�I8�������>��� ��[A�ZGg���3�bX�w��$V��J�:�,>}�ŏŕ��C��P}�W��Щ��F*]͹�%	�l{̣�ֺ�J��]��W�/��w�z����-u$���׎i�;�~b��	gu�����rHIj(�K4U�q��Q�{�MMM�_Cӻ�����ӧ(��񥾴��R�-�ۛ]����6nC���5�^`�Qy��d�x���f!U�)�۰s#�6���ţ�� ֭�-�J���!��$@�u����r�e��u\j!��4hz'�1#�,a�pQQQ�w��&w��5���	ܢx#��7�,�cO�L��	o���Q/_��̵�IŸ�ͱ�!-.>	�\���g �*�f]-��Cͺϫ��ߩ��:�����S��zb�bC�[�v�7	��!�ѩގ%��h�ie�(A�{���/���vm0"���+�7{ݗw���b6�����c�v ZI���n��sp�nLd�����i=���E#����?S&�.5�'?_�ek=�nb.DY/��?�D�8A��J �Û���mOz����ْ��a5��)h�1J�G�O��*����ݿ���%:�M0�,�A��)c>�ٱ�U�nѰ>��W��{y�-�c�R������{���fw#�U*+m��8pu0�%�A@J~� ,׬��G|n��{Z&G� RQ5���ue�H�bi诊o߀�>�t~~f�t��~�in��쇂ԁ��WZ�"�]��_	3s�?m�euu���_����Ct�JVi��2�~"��S�͐)�ܲ;��m�r�E�Vt�z�� ��
�����*b�V�^O���ܑ������ϊj�/ߚP�2�8X��#Ľ	)W��RU2U!���[L� �?�p��x-"�<<�'/��%b�Kmm>�%��+*���(��Eg�T�b�@8s�▛�s�[�|�R����\�^�
���������#Z::?�6T\*v��y���p��.�M�L����e	���M�*��fi�w�c4?⶘~��XyfN��a�E����5�����Q"�l�B�R�Ϥ�VL�}
 ��v��0Bw�q��!��c��'��f��m����v�*U�l�:0�sEr�^Bo�'�l>WQ��S��y�8�AՇwBe���x�5�/'�K�}��_nrc��m��	A� /���-�/��r�-��a��4.�_�aZ:4�T۹-8�˄�:Ku�xD^'	��2>�|Q,��&R�T c`�zt�ȝ��a=�@Wa0���-OB���RlW����"�Z3�m�D�����%������"��J	0]�T��
�]���^\� l�P���ʟ��]�ʼ%���e_������]Í�����]�xI}HL��	;X<��$H�l|�aa,�v���$7'��M[q	������5�S^38�hj�~u%Ѝ^$��}��γ���z�f�~���w�x�Qn7�XXTT=}�ex����Z��b$�����0������!��1!ީ4��o���&zyv��կ��E�#umeb��"W�%�in�Z��fC�8�%����z�Cq���+0;䶏�QP���x0u��^�>��qx��"�"Ѽ�+��-��Q����W��a>"L���}�̓w[�H����P�e�Muz�V�-����2ѐ{��`S�ҝ�����y�Hq����t Q���	q�P5&���~��PVQ�;�MOv��0�|�qP�n>t��L��K�Ta� ͭ@&���[�f&�e����\�!R|�N0��$��A�G.	A���,+)aȀ;$8$DB��*m�_r��R����!߶$��$%yc��!�k�i�ţ�
瀅ￜm]�iB/�Cp�ئ�ұ�B�Jo� ��m���h�G�-��;`ia��Z�%�v��İ4�2�W.9=���!�M�����8�*-#�t`�h��Sa��������U댉G�Wh�c��_���97$Cb?I�~%�Ҟ���:\Lă.��\v�-qZ�G���][�0 <�w2��l�\W�Ѕ�V�$Sj�J"+;A����|�;�Fh�	��߽Cux}��*1�h�j8!h��h��A]�"�������3�й)C�v�/Z3�T�֧�'���ו�	q@UQM��g��=F�����Ǟ��O��88ϝ��^Q�;��m�8&)h;-�\���Ŋ�o�d/=(L�b�Nt�+Y�}�Afe D�FER������V�dM�檴���j�曑a�Tҙ���o�(�z!��%��7��Pf���Y�#'��q`��q{�2��ˌ�r�������W�߫,�$�3��ܚYa�F�k	�� doMMQ����d}���gS@]�`k�+�S��j��)f�~|dbf��\�IG�0m�����ѝ����ʧW�]�VU�����(5�稴�/�Р54�X��CY�<;��{�K�3�׭ټ���3F�?گ�_v >���C ���>~��822�ӝ�F	�{'az�|���0�#E�N('��w&�:�<Pب=`n
׾��
WB��՘S���Q���sk�Wx�A�äU�}�;@�6��yq��߿&,�2�D�Kŏ�y̞x���Ƈ�΂�Y`V"��*�P2:*�L��^��РlR��#���c �~�֠ex{f״�pcN�]�>��xb�]a�-�S�2fff��l�l���9\��"N!�����k�R<GBzٕ��v��GW�ﵵ�a�T�?z�M#�G�f�hG�P$�9��1�m���v��\���Uº�{Ns�����v�ڸB���]��������R�h׊X�4������ 7KŬ��cʪ��5�j���:�:z��eF���{�erCS�!? �4}1���Q̒�О��~wk���7�p����ZZ��@���ա���/�^\�����,Me�uuU��i��>�e��N�V�zc�����!ZIU���������}I)I��5��bM %�}�\�m6�F"g�*��ϴ�s�~x$�L�J�&pZ/�s������/5+s"sΆ*�d}�������1t���15�{(��p��E,��O�=��ǰS#���tT)�E�߅��Io��v�N7��ļa�v-LO����s���&zUF�)F!�7���R��d����[y�UO�0SG���t���'�H&��h�M���Dz�șϩG��qT����.�_:�t~S�������_q��6KO��b�AH��n�療�
F_���a�Z2�	�� ]Y�"v���7<4�jMЏ� ���tW�J����W�^ �賴`�&�����p���Z�
l�d�k�<�.�y%��RmD�KVNv��A�
ʞ�Wo��s%�T��L��4���y���������]���'�ؾs��:��]z'�e���h����#�W!n�;�#��V�\�����2ya�C��&�ҹ}�b�����ysnՏaj��.�3���W���k�ߢЕ?���q�C<����ښoZ��[f	)9�LfӏU̱�S�!?���s�U�1�M��EM<��^�>��C<,tF����5D������c�k�	@�삿��	�����^6Rc�)/u5J���J�c"߇��	�PshP��Ό�!׭�Wg�]f�
#\d��s�0�Wi�,�O�xb }�3z�+��j݂V�݊co7�cqqQ�m���M��ΌNR�K��4�u������;<����'-'ͩ����㪛n��S��W80��jII��P����D�j�#2tjі@�/I��n�z�������e�HV"7%�C}=y�t������ڋ�(���yt���,�l����eR�ܵ&��v��
�����]�x�w�T:��E��/P�Ԡ�B���'��{�b�阘ڄ~d��
/�e�V��V(��`�Y�S�3����������W�ͪ0�ɪ8��}O��s��gkU�[Y���`��]^�°��lTG��K��P���f�L}���H��9kl�����Y��4���K�A��������[aq*$��߾bN�Ü���k�f�&B��{�cb�4�	�v�^aZɞ��Z�b�:�#XBn8j��j�Ⱦ�O�U�v瑱U��^Yybu9�ޛ2[�r��=�����-aw���e��Ê�4�������rW�6>����	S���]�!��P�3>�y`G�_���}����C�GK�r����`VJ_��@���|弢�>.�ƣ�"�C�m�\_"M�HJ���3��ǋ���袊��=ݷ�R��d'��;����ň��(QK��^9�z��F[�2�g�5'��e�_���<}`�xl}xG������O��E��V�]����[q��_��XZo ���)�S�P��Nh��Kn�����R��6O�x���N����&n��ƶ]-`􈻃�`E1	S����,�oVV�6m;˅2��ϙɞ�zt���w����Q�]X���E�QN��\�FC���P��/�7s�T(�p�x�o)�g�l����<r�\���w�>����ig�Ԗ���qWk:���g�>[?[c��+S��gw��O���J�ŚJ�y�V���8�kِ��+0	��E�g�G�ɗ/������`��??"$L� �^RA���!�-�?^�qT�?:�����Hx����v��_�~oZzQ��Ԯ�p>n(mp����uJ7߾�e{����Ur9��z��r��X�V�~ҏ�O��3�m�x�O���
�' ��pj������!�&x���V�|��
)y��bE)+��a���I�@7��s)"��/�E����ٕ�\��f�*r�)O\=�ٟ��N��s�������X���I�T���%��6�0I��A�n��3&��|�@����9e\�E���8##I&�����B����+�9��j�b����@�Aq��}v�d�j�����L|\ͭ}W�v��=ћ�����)�E��z��u�lf����9k���k�������2m9�B���#�ۯ�"�_mp�S��y̿ru-���u:���m�:��S<L����,��X�#������*�ِ&�I���|�rG���c�!!�.�j����m����Uh�hHJ��Į�uo1�>V�0p{Yu�����&�{�y��v����_�O�T�;h�7���$�f/=P����Z�H�^�&&�)5��8���3�$!bs����[��Qs���ܜt�A�EE[T*=ٳx�r�{�^>w#b�wS��7ǴM�F�`�t9�r4�=�݆IJ�n���V�WSu�K���R��"	-4�߲}�����.�W��_��&�o��n\�x��X5K��K�#�o�v�cG��(၁Jl��2��%�P��"yj*���FC=�0����<<¯���}yy�4GMF}6mʴ�!����f���г��qe�qj9��++y#N��S��U2p.��y=E���������"�n��*�@M��fU�����;|pu3�r�y!���_Qaɋ�v��-[����)�3��S4�{*���o]&�R��/b���baa�������q*�wr��qo�,��6�Ȱ�n����&�?ާ&�[�3{�װ��|�ޟ�_��_:�M� b��9_d�����^!���w/ݢ�Hh��+
˝��~�-�gK�$3�*��0�d��%&��|�'nx�H�������9��R��Nd�ր�,8��}2�x����<{f�`�Ţ�3���!tS���|�̢zz͉"�R!˺@_NΗ�7߶�����"C3oVen�P��,�	Y><�i������g��������xKssZqq/Y)a���8P���i�ο����Z�[��U�NN��~�Pc,�	�!��^tOW_���eg�K�ES�UȂ�xZ�̈�X/>*?��o��.o
b�4R�ڕ�%j���|�L{�J^�}�ր�M�F	N�ӄ��iJ�vP��qU*���W��J�!����8����"��ս��_Z�����}jy��R���������h���[���{�o��R��zr���T�M��G�dJ�|�h����7�F�K�a?�`*�!�=����q	ߡ9���6�G�J�R��-�x�(Q��ﬣT ����^DF��\��3��(6<*.���g���XsX����%+#����5� Sɘ�
�!+3�UL5��}v��������FV�<��	��Wx��I�S;2�����rv�I��%+BѧГ�j
g�.����{��+4�������X��~�� �!���k�GJM����eճU�]�$R�z�β���@e��JM4r7�4R���Q�}�bY�_D$H3���������Ȩkp��g�@9&�)>��y�bٚϽ3j�K��}h��q��ԩ�w)��|*���u�Ϙ�w�����
�@Q�"=���]�K���6}=r-�>Ѧ�c$]K�3�a{KP��ԭ)����f}���9�"B^�x���6`�����<y)��dۙV��׽Gq_�xS���YǞ�Z����şf��V�敋w�ʢ����]��GTDԔ�b��ۄm��0��j�Um�\�iU��B�z8����+�ZN-��dJV2��G1�!gDw�!�_��T��[��G�>٨�o�No�qk�sw�j�2Y(2�u�6Y��8�� N�>���Y���	E�0uz~�n�R�l�Cxt߶�Fq�Ve�b�P��������K%ڽ%i$�\�2��Y��z:~�U��0-�a�SJ�	Ǖ3������D)�1�������2{�JК��3��/}�_�zGqa���\,z��W�iB�x��"j|L���ߏ�Q���l(�{�v�ـ����߶��u�U��"MͲմL+��sgM���R��"3n����(d��#�!|z"8;<�fskk�#b�k�!M`R�s�\l�Ǵ+�,w���	{QZM0<o�X���V%
�6���b��ؙ�ke��N�&*%U���E횂e="cGa��$%�t'�-��EM��
Dp�۷�Cf���Ń�qG�Ht�4����F%`��~�2o�.0�<�ް�*�L�w�p�]yCK�ꔭF��\�m�*��A3�h ��Vh�˭���]�Ѯ��"�mzζ:�<��yʬ�fȗ�t�NR����o��qcx���P��LΔǉ�/F�gr�dk�G�o���F�	�Zx5-�{�GDxu|���g�)��/"�П��r����MF0��o�CdQ��?�0��̺0U��jS�2KQa�!�y^��Zݰ�%����,\=��R���o	�����^[��dg��L~����i��Y��=�@��Mq��c C;إ��s�/$I�-=��G�K�G8IY_�?R3�����J�ts�7#���:2䴊�����:��by�;���Ro_d�(���=q��f��֢pR��ջ���b1<��W�n)��DL�OpwSlP��=��<8�23BEHX�:oUշ�t�U.����F�p��� �����s2�#���P���;���|uď�4�2�����Ħi��+5^�#n��Ӌe�q�����ߏK�ǘ^�#yg���J�v�����OV�t+�4n�ۖ�5��F;Vk[��ߙN��B"�c�ꤘ,�=%�S	Q���KU���r�Z- ����͝V�����R�4�m���7���Wn�tƋ�L�rs�:F3�`�� �����g	��3�u�y��b�^����J��W���]�w�6�ȪҾg�EQ��|Oո��m��e�y�����.��L'��mz�BW�ݳ���o�O�U,���rq�ʭ�˘_X�����vB�?���7�H3�ђTj�O����c�8�>�%uK�Y�׏��ϛ�L�t�'����Η�nZ�q1��BV�_�:p$V9��ᑂ?0 !�5�쌤�<A������(D2{h�\�Xײ۶����+><1v6�a��1:�����i�������~�"K�A�<W¤���侫*�S� ���-;�;*��O���������y��;�]t�2P��.�ɍrr�aV�ѝde�z��/}.�)k	�n�o	����%���;��Onl�/n#�#�;h6�
�{R�^V� �Щ�������$���V~�#��Kb��s�gl#h����� �#�T�GrL&R��)�:F4�F����Jwb�]M�}��~��U���t�3��F'/^Z%���MPP��lb�������}��]�A�Sy����Gz��Toe�gļ�pT��QO~��~�F��S��&9X��\��͏v��D�[V�D�8?��t0���}���$]����ֈ��?k|�g�\-��ip�s|%B�P����G��"����TKG�&�D4�%Tl6���Jp֌+��h1�I,=�*s�%���;	K�Ǎ���Z�����f>���%z��c��;!g)%��?~BKN�Y��*�(0��Ɇ��y}V$3X�ih\��0���?XZ&t���}z�W�^P Qug�ML��
�k�j��Ir�����f�X<�W�O%������U'�Ώ��ΟJ��2?۞�f*D��~A�u�����v�c����σ����ΤC�C^��V�C��;�G䳅*S�?]}H�qA<�̟���#�P�1��KD�rR�������:̊qsӅ��8\��w+/�o=e��5�G� ���+d2y���%f�勦@�U�x��=j�g6M^�EJ:~]z�tpo^!�L؄#xQy�ȳ�}ș���_�9� ܕ�hv�&�`��`H���D��ټ�@-��UQ�ꅵ$e�����b$FPǇۛ��G*�n]��f�`7&T]����Ny�#&�;�6m���ޕ����*\��c��A�����ӑW��@�#x�j�Y�#��}�;M<��~PQQm�
-϶��*�P������-�ڥ6��i��?@
�=\���X��^�;�˗��:��L��#nI-]�~��T��n�W���4��ύWԙ�mKJI�O��S=9��t�T���Y�W�m3�{R=�^�Y�Fv������PN�@Ӓ�%r��A �ۖy�V�#]X}X�-a$Y)H�ג�f܏���/�W��d%rԢ�Lb9��<}Ns������~�|=�ޱL�ny!F/�so���.QQ;�R����2u_bc�Y� �k@���<��Xh�t�v�;X,�{NֽK����n����g1u�%�u[�m������;���Hی��P�����	iK;S��@`�M[�Tn�%ՖVW)��L #���ą�ͭX�OYT�;q�f�H�S�q���xM�9e#�/�<�ɍ�ܤk)�-�n������?��n��4
l�0ӣ�7�\"�VLi'��f�������p���2/�|�	pD�,�-$���rz���������	����C#��N5O9�����ŋ-M ��6l��Kyr%�_Jҗ�{ ҅��p3�=���i�*V�tp�T����ó��Go�]&S�2u5�(7����=p�0��\��b�n��]�r�8�a1���;;;�:P� W���P����:'�CO-�|�p�j?��A�F�(n�b����Qj=�#.?c1g�"�5��������}��a6��"�$�^;X��tx�<�]ȵ1�:D�ܾ�?{��se�>~�GN�'�Z�"=�����f/��$ކ�8uʙ���l��ń��=��Ѣ���>Kܮ�c��	 hŎj�������ָ\��M�w�'c���C���`��SS��wj�����#5bN�:�v��?��ٻ3��` �A��=�L��Ϡ�$%Z��ĿG��n�=Q&+�Q���a��8���?�X�������M }���Z���>�pc#�<a {����^v9E�./ߎ,.��qV#ƺ�nf��	�SS�>��ޣ��6	6`=ֆt�IN~���	@׌�ĺ���J��V�g���/�c�I�� ǡ�o\:�'z��3`��`[~s �)�}]��?�����;Z��pY���W�itLE�a3��jV��O���dk��O��0���/���R*��euQ����~y3`# ��� �g�D�~�p��Ġ�_ۮЎ��n����BYJ}�"�C�u�am�z���^�c��<������͛����&^9��۞�����ɤ7(TH[A�P^}J|��\M�
����<���_]yʭ�����b��n�`����+����S@h��ܬ/���-.f�|��?�aE�'��;��m )I^�%˺��X�:�\+[�s��<v�a�������uKd&+=�-"aT���5X*�ͥ%�(oqe���p���~�1�J�v�d�.�Bj�	e�9q�rv}z������9�tt�̎({��׀��k��ϧ�RRg��W�l�����������"Y���Qw=˪�S33�ꐟ`�8�j
%z�u�O)�>4]9�Q����ؔ�5��F��c_�\��R���2�-�?�l�(ҧ��gT�8C;��7��Ψ��ŭ��D�c��u��t=�5�]�*2�ou�����s���8Y"�NQ�˶����1=�l$�x	U�Dc{��\���4Sss�T���9&-��4t�}q����� +v�"��(�i7[lR��	ao���,>¼ɣJ*�v�sD�\M޵{�P�ol�u]�ü%����G�O��&�͜���z�ʨ�\Ͷ�؈��J�s*��^�燫������²�קc;�u�=���-5h�"bb)m�P[Ys�X�^ܤ<���2����n��GNN�̼M�wQ�N��hw/���BY��mUU�z���5>Q#bX��xa�>�Z4������5� ���Vs7��&�����1-ՒCHӆ��Y����<c�=���d���U��.o��t�򳀡*CM���6�.��0ƒ�De���'y��7�p[��a������*��'��MF������"�֢u�ȸf�iz9]����6/F�۸x�~�po����$%|%�����=f�rs��/evR��0����N��koq���3��>�G���ս��B�L69 #��ΞL�39abQ��充(�Ĉ�"L�Y1��`�؁Bn�Q�h�OG��I8�Ƈ|P���[�U |�.�Q1ѵ�96�ʩ�*߉�[��` HdR�ӶK)6��]�G�\G�-��$|��6���qoN�6M���s~n�9g�e��댻�>�N�����\S�~ �4R���h�qf��1n��{����쒋"�	G��
 ��؇��k��B��d�S� � E����@�<{���!2%�ڃ%��*��2>>V�Q�-n��r����K�[k��1j��+�?VCR�S+���;=Z�X�a~ܾ��߃�n{I�W���JԹ�?)Rؗ��]%E�ˊ�F�K��G�U���p@i�&0�$�(ڀ���\�H�e�~��;�S#:E�{y6��ݹSl1��_`���E�"��"U�:�����Z`Ԓ����l%Cn�����Pf�!�|�fƏ��1}�z����!�R�
�\��#�����	DT��:�3�)�z������V]P��]�����n�3��c�9\�r�Е#���c��t��w��x/ɧc��(۔F��vZ\S�o�������ԭ`A�qD�N�y�e�.�|0_+�u�S$}U�oun1/��'�F�?�^G:�����]�颰|���8��~��%6S�"a�ئ��'..��f���(AǟNAI��?B����&*��,�6���;͖߫_���<?���
�F��\��Q-���w���f���>=6��Cki��X�Pkj�_趼}���=͔��jU�x�1C�*�2Af�"��/��hK�	�5�����^Fz�S��6�k�l}^����z��΂��D�ݨ {W���������ܾ����VR��(s"2���)�<e��G�
ɔ�d���K��8d�y:�y������������������Z{?{e<N�7y��c�g���]�p��{��a�F4"��G���s�z,��e^���--I�	�qR93]9`��Ʌ>�T.£�Q=�u3tƉ���O?����+�M/�B���u-�qz@_����+�Y��b�h���*�W1H��Z�J�K��Q$�Uh�PS����/w����� (Sop��3��=��Ӗ�6��s���e ���7�[�Е� �"��!̎S++u�b�;�Ф�w��vM��l�����;?�ʷb�"�
��>16�ȡ���H���x�M�|=> ��U=ɮ�bW��h�#���=u�q�o�ъ6�Ϻr$�
�ښ�>]_G�VN��%I����W���iwN���>��?��lEҙ���\�	��s�-�9���T͉��*�G��UY��j��	?��o�v�y��K���X6\���J===�2�x��̰��xNCGG]lB�B`]lxb�f�m`%�u2 s�u��#�$Td��j�@��[�3��OB��k{���CC����M�ĩ��#�������յ5S77-`~-cJ�⭏J���������im��O�I"�otn�+��^mn�x'���d]��ӨHE�i\z��ħ��ka�q=��W�Sv�S�������~Zoe$����ϑj���y��E|�9�C6�l�<��\��ۆ���n$ջ�
@�������U�����>'��T�5�JF�t2�D#���t{���Z�q<g`�ূoﺒJ��^��8�Q�]m�� P3�4��Y�kz��!o����l<Q��E_�1c���%�fTj�$Yz�(��G��uRYf=���6�=fk"�nД?dIS�kvnw}� e��b\oڜ��ߎSq[G|ο�tɞ���A�j��$��x��r���\���s]9��&��x���\��(Ca�wd���*0?�'��Z�f��eJ��y�*��rh�*O�f��x��&w_�;Q�Q��/t�~Q ��c������r��!/��+ ��p����3�²Yw����s�����ޤ\��ؤ�����+IG\%�u�؜'Hs����|��[�ɕt���j��εZ!+��	�a]E���t{�O9��AN�*~����}�rt�9S�ӴK0��B��~���@f|d���,�=M�36[־S�������(�2O���_O���4s�������L�fs�YDr�X���5��=�-��aڿ���h���Ŀ�rd������ͬ|��R��vo���X��� �G���5�'�k70����	������6x�MR�?�3�	оzl�r��d8����+s����k���Qv�������_1�Տ٤�,�~�4U��ro������ʑ�-1�zc����E���|����_Q%Λ��m@������J�%�|�)H�G���Jp�Dc` �N����%�8ޮ(E ��� �œ��t�S�l��%�*.�Ո����^T��|ܯzcN�-��S*�Yް��Wy\d�b��ɗ�׾333s���I8�z�Y�@ *����v��y��IU�rkӼ6?G��L��לPHQ��̙I��pk)��1C;ٝ�kN?s��-<a���8%����5<e;⃿>ϥjcs��<'M�k��1��r�t�F��o��Bp��������m�j��zC���y�2s��G|��s���W^&^�|�uDu_Ky��oi ��R�:��w��		!���a�Pu��n�m6�m�@�C��/�^9��#������w�4<ɂ��T�j>7��d���[b�&(���[�{"N���gx��29���ڕ�� ������<�-at�����.J���H��+U�n�S[��a�R�@��6b���
锷<.�kd/�n�N�Qޮe�������Ӹ�Tp��s#TU`ֵRà{$�A�yڪ����'�T%������K�V�$H2��țm&����ܘ��m�\OO��W�%�8m��E΢���\h�)��ɼ޾�f�P�?ldW��l@���ت<I��el�a*�4f&��T�.�0M���a��N*$�T�B��]"ס%��3���"�pϪr�P�5�S3��F��຺�1ן�c-�Y-�A4�lܓ�L�y8�R�#�o����c���/���])�ܽoY�
T�w:?76�vquH�jƛ�4��x7^_�����B���`�����w9C�\fx"f��ڌt�$3ol�붾�A<�	ao�W{���y\{Gl���0�}��`q֢��C�!�VIvw��5QXª7ķ���y��''�g}Ĝ��w�5|Du��#��lmm�6���*�ԕL�#4�Gܓ��L��Y`A�g��ͻP��P�i���c���i��Xf�$.���Owp��NZ	7Il�NP�M�w.RM�N��;��6�!��&jcc���Cb�	.�����C8ĶRU.�c�����L��ӛ�Q�.��d��SWӾ;Zo�m�� ���$�5���ͫ�Iz��YT�N�&yR��K_�Ϩ�(j���*�����q�q*���MQ� K��pE��$1��GO�8q�<��JkF���ɘ�����S��R��J@���Q��ۋ��Ɂ4Eh���Zuu5y����4�g��s�u�����֓��>`!�s�-���D5y�W�'-�����4�����q��u������G8v�m�L���U�m�&-S�	V��]V	��ֿ'�I�h�nnk���B�DF^��eQ��aC�@x�I��w��p�ǿ��� �qVȾ��E�Q$����ׁ)O.�<�'��FR����c����b�]_md�C���#�2AhoO,p����i;	0Ŷ}��os���b����6�Fܩ��v��8����\J���C8�u(Bg��%����Y�fD�@�!��J���wjKKޛ�BJLҟ���pWڵ���Ԇ��hL'%�[<����}�����(�j�3��=|)��S�Ƨ�N����r�D���J��$
U����Q��ֳ�n<X1�q��k)�ұ�	E�+M{�3V��(lE-�3i�8V���z���RsЫ�R����b:d6�B2dv�|g�K	ŇTE+�W�nFc�Mn�[�0s�� �.2��`�	���a-�n�:1M$vv�pr�x@P�kPU&W��5E�TxǍK���W��3��e��0"|a=�x���{GR�IZd��]9R����t1j�is��79j����p^m��h�y�lgC��Z���B�0N~8ም�ʃ8��}^���lҗ��89��n��������<��Qǹ���s��K�{��޶La�ɤ�����6]mf8�� ����������Xmq�T���::�Ars�D郣���q�����)ıi.��jK�V�����Z�U�P]I�5��;8���q��r�I�Y�&fY�/�.Ǝ8�d��3����Ψ+G�za�N`c��RR�"�6�uO���ﮇ�LP���5IcT��3�'�ɤ�s���:�:F2j��h	pM�k�I�]!�B�&��5������чT�!E��$br;�'��>+�l4!�����5�7����������W��K��1���s=�S��.}
yF)� ��ύ�DR.��D"CXrk�<<ԑz���9���A+�]v�mo�Ӑ���+qǐB��YW6��c�������Hȹmsy⚨(g�q�[䦴��!���4i��]&���������������>�hOW���?�(�ȝ�L�_$Ĭ��]΋�WJ���u3:y�1EU�џJG!��~(A�zn��?��������?8�[�O)g�"*M�넋���� P��u�
���E:��[X���̐����v��`�����S�yn�����K:u}�u�ĉ������!��.%�LYynG���V(����E��>�����g
+,�7�6%��{/���(L}�F`��"��@Jr����BM��'�	И 4��똥��=����6zN�j�t��G����ROҶ+9
���-`(��l`���M�o�d��Wvek�ܿ��;҅�&ѿ�R
E�$�Ǐs�|O�� g<TymCk�~��h�x=�|�ۣ���F-�̴�K��g�+��T���i��ݕNʽAT+�B91�픍ا"��^�`��%��Pz��������}m�uL�$�RAtc?����C��%G`jYղ z��Io��F�^�7\�2�m��KI�ZNRjK�\79ٖX?�w�oe^��-��q��4��[�E<U��k��t���Ȏ��O�$YJ�'���Ki'��\���)�P\�㋒/�@IeF��nlFFGw����u\P!QɄ�c�e���E����#w�K�,&��O�$l��3���S)�r�"�X0��Y��E,���.sz ���>��gkn�����4wx]�ݍ$�v��CR�'Z2
�VWW�f�}E���O����Ji�X �[���XH��WE���������1wY
� �+!?7w=0B��=�Í��� ��հ�G�J�EjP��-�L������ԓk��y��g�2a?��w�m���+қ���A�cue%UiH�B��3?�K�0'�E��Ѫ� A�d�(E�L����qu����j�����q��GU�Ķ�c�1L�&�F_s�|>�+���k�륃�ԟ!	7�Kyyy0���b��)�F��燻�nȩ�;��q���n��ſzz��_Kc��ݥ�|3�{#9��چ�O��x�r�f�[�����B���ȎK[�B�>8y 4�/WL�y� w5wc~}&�v~U�z�8�[s#��Ɖe�خ��PiaW����4P����7:j��$X&/e�q�����3iO���{#n]��Mv��+��2�D����֘��n=S��P���`�B�$#�����wE��`U�P8����vc���M�I�Pe~EK���5\���M�+n�s{���7�n1�2a���A��)0EAd��qp�b/�pɃ,�z/�e�X(��b�����"BA2*�
�Ɓ��.��9#x\�}�&l�r����:�c3�)Ux�`�߾�zr��aTR4�L������2g[VϝEH5ZA(��Qos���k������O+K�p�����M\㊖@+�)��������P7�bZ$��+�9���ŝ���4T�aȝ�%F��	��Ϋ���LQ�w�>��R�@��0?���(�����_�5��K�IS���.�	�ek�K�K�����@%�"��������iy�]�.�(�=��6s�	�'��2��Č�=c����W>�"?��,�=3wj��9�v�X��˿��-�u�޽C%M޻�ݭ\����kvc��p���p�h�"-�)	�n�k�s��0��|i{(�z6��Łf`W��_../k�$��� Ή����p��Q�{����2��.+c*-��g2���I�0��75��`�:�X�Kc�W'���qB����S�^+E��<��L��r`����Z����UQ�{�����w����� O&Ɂ)�\�j�YI����v��rݨ��<���⭽�6g7'�U/�ٕ�YM��3�lv�8�?���}�����.3�r�Q�|a*�Ag���ؐ�>n�����슁�5Zo�.��8J���x�) ��'OI$�WT<��.�=�L�S�@�ԉ]�`Ӿ)k�;q�<�<
���w��ԏ$�d_����J�l�]� �]hmlֿ�1�oJ�<�I �f�<�>!S���u��*�{����/͌��<G��VS�s�1�j~}?��M�7�^k���ZϝZ�Q���<�l�
P�ծ��(oڡ%2�Y�6mG���?W�,5lF]��2�Ǿ����p����o�1S�5?s����Q��+;�7e7_�m����d�Fv��o�9���{����}���j��v����K�[�"��?��y�;���["Ҥ]�t#֬I������h�[s�a���3��R�0�Y���,�o�yCai�C������Z���+4�]�� ��g>�{�7�$l���IK�����L��CY�Sٕ8���#.��|�\D��&�^d����z�"�Pk�es�wֶNa.�+6�Vz���@���������0�����p�'њ9�K�;�`J!��3)�����*�-�q<����	}�$ ��`SS�@��m�'���z�i�w7�VB��N>�&��l��Ý?�U�|�N����>�λ�]��{@�5�B�ҫ�2���Z�Ql��{�Pac��\�?��^�7;�O3��ڰ�Тo���B���7K��L٫�u���c��sL��2�
������o�nv�j}˾�D��â�z�xP���3�}�����5 ��B�;�-�����in�!��V�4f�_�]�JP�Q��uVB��0�7zGW�Uߔ4�I#�����R��ja�;-����^�Rdu�^�e��j��ch~}�=J��]a�ô�vH�'�I�Id+
�A[O�Ʋs��W��gm��'/䔯i
YD�Ƌ`���3�}������C+E�AQAOc���z�sY~n��8��o�l�Ɋ�Ab;�M�l��w��*O����&Oj��*����Ed�1b�Td��`��AB�A����\�i�|Ը�G�+����s���|��/}?�)ģOtB�:e�'oo�r�ӡG��~��9^T�y�1H,�C�p�Eo!f��h���))��߃���L�Swg����Օ���hq��sv��x<��z�3���������U�oW��mr뫰������gZ].U� �X� )�ֈ˰;9x�
�����mG��K�Lq�Ys���k���E���;6��]�z�8�{�dʏo�Έ�O�Ʒ����L���8i4�Ŷ�_tk.��S��v��o���o�y	��1�"�3���E�Y�o�{���c9��Y�r���y�-^Y�w����]R�\U�����Z��ST�����=8����-A3�{W��ɲ�{�r�m��hsc$�c�s���� D�x��jU����}�s#�������0d�Y0��|t,���_�$( ve66;E$� �wm���$����O)D�*�*�SW�����:_���\������P��ݤ��J"��Chͷ�fw6� �è�b��U��z#ǹ�j�Y���`7?؊Dy��Y(�S� Yûo;����Sn!ݨ���/Z9�����^t�b�s�a<��)X� S��mos�yw�`���B:��sc%�j�'v��uW��h:O%���<F�����z���h�5�!Ѻ�=M�UxpO[�%l���i�6O�z*J�es�{pn�}Eq�;˾�[9
W�>:z#����j��W��8��0M����.���MD�;Ш��'��^�Ċ���"�p/��ϴ��P�b����<�U����:�Y~h�O����1b�����\��Q���� �7*�|n��F�˰_%V�n�T^�w���v���Cv�T�*W:_Iz����@�o �q��ຆ�����y����"�ЅR�V\TH��{���9ƪ�>oV��s�r�Ү���X�_�yh7��TWË�6,����	�+ͽZ%_�n��q(�j���
w��_�7������J�g7�=���R�?M�6�+,YKG4����"�]��o�V��	��P艖����!�����ݑ�B��7�Bt�RP���e�r�@��dٵ5���iش%�u}��V�c��c��K�l'�)D?hzU����W���u��C4=�16�یy ���x]�H d�<���t��l
�0�#5D{�8�b]��~U���#*o���ZB�t�׎�/[�ʧ�Kj�7�����cR�mnX�!WW����_���u �|����>���'�����ʴ��q�ܯ�T��#@�ˊ�ѻ/WrNC��~�=�B�`TS��y/��*��b��G�=��xaBl;@��1ԙ�d�`_���u��1��zS�^ʍ�S�������� ?e�}F�^Q/��{��Cþ�F��P3� \e��R$��ޞܒƅ�����u/��*��	v�� �IS��u�A��X��	 ���� ��X����B������Z��彟��<Ab\mƣ5��R��R�WiT"u,�������%(_��h�zǳ&�zS���|��0:+
���Ic`o��.U02N^���3!C�`�T�n�ʯ�2�T���m�܄<�s߂\��,b����jσ���-]\D!лFd�k:�K�C[E
���|uUr�BQ�c�r5�ޕ���O�ʃ�&3���ނ*k��j�,h�:�Fj��R�!iX�@H{�gw��W���d*�lg�	NjҮ�CrY�i*)A�XY[�OC
2'W���q�_x �p Vy�jZh�>�uv9l�dP�P/	(���u���t0#a�A#v���.�� 2EK�;xtYL�2��" ˢAx5�\e�e=���b:)�\3o�.��:�4>7����p�Cg�\WVO����BM�� ��uec0�,Zkg�Zh6��̰r������P'Z�eL%��[�Fr%�jo/��ބ}����0׋�zT*���Xg~��AI�ڞi2c�V�RLP�-��@����G��SZ%v�|���/�W�H)3n��(5vJF��p��kl�K��e�m`<�lR`�'*�_
 �W��L��=��,����L��Vv�'�l�>d�d<��=O@�q8�*Qx���\�W���( �=)0��e�!�Kn�����5^�=��z�'��+W�=l�5X��R�Wh�eO�s�U$3�r�F���h��c�! ��u��ϛ,P*�6�Hd�!t�j����:�Z��d>�&؀t,���+􊀀 ~Lw�D;����Z���G?�^P8s�|*�
\���
�d�&7~�G�t+ܷ?��t���Ds����E�^����H�.h�b+�,7,훖eK#������0d����Q���0����>��aO�#��$p�IJw�,&�\OD�n��-���[Bc��܆ج�)�x����+M�s�,�R�4��9��f{�ZJ�M
���$��a_@�a��;h{�$Y4��� p��NҨ�z{��X�/�br�L��ˁ��\��?�W@^��mGq��l�E�1�r��7�a�J����h�����`ߖ��m�}>���U���a�վ2g�ܷ�̩c^{(�	s��]�O��}=E�s�E|X����u�a�l��W���Ѻ���+�ڠj��Q�̝��
3`���	#F����'�JR�4�O�:I���T�q�\�i-�R{��0
�`���/��ױ���͉8J591����Ϫ�P5���0�'U,"Q���!iw�~��l�Z�~>�t2?���z.Z_���+���
���͂h_d�&,�D���Ǌ����`=l��K�at��^��u����3�X�w�+¼�yɟ
PO(��� ���^m�B,�&3䳩���)�����d�`]��*�AXm�J�Z�!��c�%�?��+Q�sܯɛ�
����?�����5GG��/�K�����`UrƲD�^�w�(_#�Hu����.ps2s�0a
k���l��+T�"T�K��9�lb���2�tI���٘��ɺ11��{ 5ہ� ȣ�{�_��z����#g��y�+��{�U-\x�_,<�q��a�>�k��Т*r�v	L�;�������#ǆKR�|�cj, �]Ǹ�An?���"��8�����Ue���Y�]k^T���R�)��Q�OA�M�*V�� �'ݠc��:_��`9X��aI��r?�������l��(367:�����B����}2\3� 8ޫbbb�Wr�
Jp��B�����ZQ�4ܾkY��g^���<�ʤ9z�9����i��-R.}WB��4˜�L�p�0�t����Nj@�g��"��q�g�.�5x�A߽���V)�y꭬��9�&5=����g��TЅ�v����Qn��Ķ0M�,ڧ��a�tÁ�s�WSZ�ͻ��&�l�CE�����x;"��R��R�D-�d�i��Hl�
�2�j�9HI�������U��̗T�(w��j���L����ۜ�9'�.���?��Jm=��D@�vD��n��a*YZ�#Q��VUL�a(������n*�X�	�j���׬ڝB���P���5�z�X`r��C�{i��F��j�������.uHBݤ&������zxbk���.t�F�ź ��=T+��Q���6����9@b�7���o�L��m�s���Ֆ�0oMceMo���f4N.O���� %lV � ̂�^�j�$��PX��ߖ9���d.�S�e١!˧L�@ޱ�]�����d��N�쬹�$u�	U��h�le�~i6ܧ�)0�Y�&�/Tڨ���h�ƆSs������ZJ�p�h�rL$T��*6
Sv�م��:E���tY�@r5,�,��?���e>��iQH�j�j�;�o�$("�8�.LI�8�[���o���ؘ������c<}�k�R�X�cF�'&�w��S���!v^b{�F���E�Q�76y(��T�?[z8csa�N���w���d�"����N�TC2�A���v�A����Kc�z� �~F�ŋp�`m�������ܧ���\�Y��1 G ߪ�A:-b3z�c���\�4d�cWC�7�]�5��/��N�HEf�kp)�a�}v�T���P�"Z�a+�!�i[����}]E~B6�v,��>��)F_�sL�X�g�EbcU�NH�U����m �zY=�������F��5��X;uq;wa6�X��+��0@�2OK$�v�D7h4 F��v-7��5
������%�sw&M��_�Z��4�,4$  x�C��]�� ���0u���
h�a�ps�ѓVi���2K���TѠ-�ݾ��Z���m�k�Lx�jŬ�&�}ժ���� �;�j��\*���ɲQ�Us��K9�|��x�gM ۞}l;�:R8Ar!��=\Xj�kѵ���JQm������ƴ�]1�]�a_��E���5�}x�x�\#U��!�n�-��\���� Qҗ�o�m��L���24F�[��٤p*n_�������Z�Y],2�*���'--6���8��0�֣������+��W�>K���������� �WG����2w�m �Â��[�e�g_a�A
�C�8�����4(�S��XZ��%#�5#@OX �dr U��Rvu*�&�bol��)Uᒭ(ޘ(Y/\���4�ZW|�ysNI��LN�2)s������n��3�S����::��+B��sc�==X��!���� ���pc�ԅ�>�V��0ƳC�=��m��`�0-}�ڮ�����w���rnl�rO�I��{�o�����t^���0���7�����S_�/e:�ޑ$�U���ӄ�!/J0���>w����h���Q�$�7��4H�ŎI7�R>�AE�_g�ߨ�/��k�nZ@.o�b�;=�O�����ɓ�20��c�	��
��(��_�(�̛ï����Y콇Mщ�S���ׄ�#�Y>5�$<�27���%�Kl ��R�dx�]d���z������;���?��+Ĉ�����ϰ82әU��S��GxK��jd��W��Mm�W��H���}�]_7$e~p�6�M1�ٖoR~ZQd�;*3��<�R��]k����l�!�ڡ^xJ.P~�X4����
�`vؗ7I* ���� ��I��9�2'~ϝZ�hl����;tLL(�rC��WRH���IP�<�a�k�N�����b��ls`������~w���|8��B��PDj�����L��P��ճ��@��8rG#��q-�m��J���i��f��$1�w'�@ŭ
������,�)�EX|let �pl��4A��|>g�}�ԫ�؁�i9P���/8
[[����\�Jn�c{�dz��g2�ڕ�u�􁳯���i��^ ~fٜ@)���=چ�12�`�F%�0�8engg�w����?��fI埁U��!2��"�F��P�X ed��|�v�@�E��{iy�q�r�H�\�ٛ���Z�W�tT%l5����{g�c`Z}l��/@Ԓ�+�Uʗ驜ͱ����1��>��`�'bA��\,���u�	.b��V��F7YFFe��V��vI��p�#����^$]Q�1��ܐ����:�)���ѹ������+�r��u�>:��o�e���F�&!�%���do���X�'�W�.+� &�屲���`����c����{����u۰���p�?(������1�y��|�3�f�X�ƕ���7�����u+c�8��Ad"c����
$�7}���x�ZՍ�ݵ^ȂbY��bNŖ����R��5��+�!�ȘJ������
|.��Q T�m� ��z����^5�a/�EP��x�Y����{�a�����H��X�Z���At��`��yXB�G�2��/�r������� 5��X~�+���=C�(�J��l�ǁϵHW��D@��.<k5V+�t@*����"� a�x�7����j�.��k��<qs�q��Bm'�n3̄��!��. �4�ѫ�G�/ʴ�*zIFE�~���諺�ђ�=/�RvPH*�D�Ӽ-9g�x��ǗJ��62�̪ڍ���n�K��»@�U��#l�w��3��.�IL�� N�R��!zg��JaH���0����%��\��"� !�|q���"3��̐׺����vm�{v���ڇ������ՙ3,,4�2�y@;˱qa� c��U�R���{� �*щ�@��jZ�9XM**���EZ(�snN�����.���7>���@�s5��͂X�V]�UG��D�n��9����9��p1�Ȇ��3r�J���7���o��?H ��uerJ
ܵL������u`��G��$��� �eZTC%{� L�>���
��q��^��>++�(j�9�v���O�j�(
9*u���6p��%44U=�5�Y�4,�˕�������k{u��
�����Y�櫋ث��9�R(�n-I[)VDG6}����T�(�=���+X+Mt�l.�U� 8`f6�m�������]x

��������2Stx� w�3�<=�ֽ��b6�%@��������{H�B���ܪI����ؽ�3��	��->�(�l���i�ܑ�����rX���r�J�W��Cfd�=��V.u�DT�fck!d�/W�O;��M�=34����s��C�)R`�$�S�)\%?"V`�yw���#�mo�(	���)^u8��t��<Ivd��k�}S�^S�c������t%���:��K|e���.�&hV���F��x�̐N�f�&�:��p�w��U�8��665Q�z���t+��yD�N�_k��A_lO��7���>��<�ý|Lk����hD��r��N����F�������$䠁�.�6�54d�̽R.��)r U���og��M��m�u�E=_<HS�o�Co"�C��K�N���]O�!NU�����|U��
�P/��K�݀gC���s�����K��
;�B��X�����3L?���1�b�1�[yJ�c�ݑ_(V��qV��LD���ǵ�\h�Yl~�ipC]t#�W�Q U�����ezL�c�VZ��|��L
������#�3/ђ� ����8�D�dԋ�ׄ�~�S��Ml�����N��]�+��4�j�vF�`q�X���I{�_'/f?�V�Ț�'5��L��t=��y�1�����=ԍ_$���\_�S��ޤn�S�X�-�J�&ƹ�	z���F��� ���"�f��9�:���z���6�g�gT��<��G]���!�u;�Ѭ�C�cZ�JvHLxZO�[��Lc�0�G�8�#��5�X6�t�FFTd�g�����[�+鷬2�N�C�����^�49�ϻ6Օ9-����Է��
D�:�����qG�g�H<�B~�|\�ڈo�Z�](����}�����o:�-Y�f�+��?>z�u(u^�ܡ��F-�FF����W�*���at_׮2I��5�#RkVI�����m3����b��q���kV� �]Ʉ�5��������ѝ����ڑ8���+��}H��f$5t�Uʃ��R�GG>�
^��������k����Q���y���|6�>?��^�Jg��N�e�vy��U^^ޟ֚q]��a�Y�r�J�����]�l������ͻ��T�n��흴�$���WEb蜛��_h��ϙ��N�������7v��n��

蹸����Թ|�[E7T�?M��q]ٯ�?\l;�~�^�n���K����<9�l,�'�J6��0M�k�:�l��*���"
e-�&���f�N`>�ظ;�-[���������&��@� �+^^�B��!Aޮ~��mk��딤����N����R�З*w�[ry�#�H�p~�wu?�k�;G��k�������=H��LN1V�O���Sa�ǘg�b�]�5�4y�>M:mV�}��yg�]i��vA(���d`���r�A����I��`ߏHm<��<CTXq)�Mى�_v{!��df��&�Xp�!�1b7A�^��:�Ġ&f^���	������G�~�R�g|���Và���������u11��O�N���9x+��JS���m�����.�,���x(�WVΰ Խ�Y#��߬��҄��_q-��]\9`Bl��ކ�V��#����Tt(��z�vB�����[Lu�R�h���=��&[��5��oX��3��澕A����m�o��]-�;�$�m��h �T�e���O
2��h�΄�x��N����0Fs�ܽ�%�����)J!�����Ծ8�2!�n���z����j�t��Ш��6Re�Oj<�8]d5x
.��1xN�mY)Ne��=k�=��$�C����,���R��^���U�夵r�˶]5��+��!i���|�<L�J����,zZs*������I;����^��6t���k��Ex����u��aM
�帽F���S='���Mh��i^K��|wku��@r��m{��R���7x�<��ᇑ��Hv]ur�8b��� �9vM�oc."�ϻ��r�+z�M'�O}I�H~�$5X���ν=n�莜K��\��U�cJr*����ck��L��]����{�i�Xd:M�n6�a<���D�N�ӟ �1��@�D�;�_�`������;ooi����|������Z�'������m����I<z
*�i�[#�/�;��3]9�9^��Ges6�foR���/�;a�j}~0~� �|�u��l�
�u8��fa-��K�^�d���n~�G��*D���v�>
�ww��x�^�>�}�U��z��oܲ���UӰǒ����ıh��9��[Y�f��}Ȏ�ә&9���V ]��ϴ�$<�zEF�Ϟ?�/,*:�0�����c������.�E=d#���!�կ�t%v�KW/��fw4 ѽ�d�hX��g`ii���>_k����Q�ڡ�E^^� ������� iɓ��5�w�_�ɖ�oBIT�B��<�����d&�|�cs�1���WL�iq��`T�� ûr�o� �S�f։n���q$[�[�T�`b�4eU�8���exX��fn�)����W�$s��kv��}"}}}Z�c /�G�n%����]YX\���㴲B�������KF�|�����:�>7cLe������z�T�$��-=��uݲ��O����v%�!)�R����-��|����0������A�T��j9��=�^0T%�/�]��Yl����x��
I��!wbw�Q^y9�u4�,�Kd{�Io����Ukf������,� g�������S�$X�D���Xs�H$� ��)P��R�J�rs������$�Ķ!���82�_f<O�<�FD5�-�*�A��άv�i&qʦ��l�4�m�CCC�?'^;w�Lz�Dk�G�כ�49���Mgdɋ6ga@?V������8��+=�C��C��� X$Xv!-x`\3�Y`�����b-�=����A�Ut����L�d.@�!�7��~�sei��Z� ذ遝�]of)@?"��0�-s�P؁�v9�r��ު�����\�%N*P-�~A�- �Z��|�_q�v*�yxq�1�b�2��a��<��Df}��ߔǩH"�J�=Eq�� +�����㊠�B��d)ϳԨ����|�z\����vI���C�y�'\��)�\|�&�\l�r���ؤCiP�	�5���<�� �� �F0tM�i괼�
�!�/��a�p�!�����;�(f��q���=��Z����`P��D+���~��<3Ҧ�Iy�E�9fS[[�,���q뷑�;��T�j���W�<�Mk�I�ߠJ��D�������o���`�
$j33�< ]�H�����Ed�����Ƣ��|(b��}Y�1��}�n���r�����1�U��&&�))�!P�}��!9d!ɘu�����;���
�JY�U:���̑�MzE���\4^(�T=���k+\R��s��o�8���؞+�mZb4����NЏ��dʡV�N�C���=��p�A� l*���H��u9�{s�`_^N��L䶞P���YЁ�q���Y����u��I!�[�����Y��X²mFF���&�g@*� U���R�5X���p���3��/^z�o%Ѻ��z�p+�����!A6��8-�O���UN�>&�$�Ա���?eP� s�}4�U�����Xe���ݯ�S���e���k��!��Y?w�>���˗�<@����ص��G�W��M�d�xir�&�k����AY�YY�c�A��bFv�����$��j'@.�Eh����5~�6VYg�U
����9m3��eO��Ui������1����������c7���=��N <aOI���U��8\�
��&H�:C��C͕�jKD�i��PC��Ǜ��7���	��֋ɦI�zMk-S���_��Ĥ��t�'{P�)�X1��䑌��giv�<��BZv3�Y��r���ȥPL��]��oX��F����a&���>�g>�$7=�@�eH���V�~��``�(5����������h���nW�.wɘ�~N��H��Ü�W�EV���Z�"�ߙ	�̆e�/eҰ*�<G�n�R��ڕ�kjj��r�f�6�t��Sb�J�L:�\z�X��[���DCW7���R�GC_�=v��m���l�4�%2��C�`���bM^a�)}7���R��ĐK��x�M�yT�SSS��N�Dۧ�yٰ�A6)G��	�_��ی(//�~�XWW�@ZsC�y��Е�yt��,~�u8��0K~�R�����gaaq�G��5��Y�����p᱒�:��ѥ�;c||9�M�HL)��u�g)ש�l��JDg�p�ȇ�557fq��.�uVr�#�>ş� ._?ޖ}oLw�"��L�{��d�Rڰ�պ����KLJ@J�Ψu��Ȳ�e�����['W��/�'��0#�2�ةf1� 2ǦnN�']"�p]�&�xaρ�I_6��v~с'F������@\W��]�x;T����r,I6��kե�	���{�U9�"-U��Ǯ7>��?�^ث��R�7�}}��9O]��2�F
C}�q�_,��m��s�xY@jo�`gwp��uX����8�VPP���yE�5��6z�,�a38�F~��U��dU���W����~ٳ�ư)�s��D����P���
����ۡ������>�2�M�������,^~	@`��^���% n�v��X	j�~�r7k;�1�w��=��Ί`�M6�(+��c���}�y��-<�ˏ*=A �ۑ�4B����'`n��/@�Nf�.�8�_�x<~c4BK�%�,A�f�NS�c@�n�Q�$��q�
�z�����,�HQfY� eAd/jC5�5+�J��m}
�u�e�:�_�k���DW"RO�w)o�Ha'�}���� Z��]"454�8�S�^Y1 E%T��B�;t��N
rk������؁9�iqbz��W�:ڷY�o�򿅍��W ��B8[Y\����A��~���4���r: �P��8R���;�E��:�fINex�7x�lvF��`���(�K #��ɡ,Kw�9^�cExU��3�;p2������ޔ��c���'x��_�ߥ�4pN��e��H R����F��,��K(�ث[8�k�LsxӚ�8��^����$���W&���H\��<y���Z�1���Jd�1G�`��ʊo��	l-�s��Ƿe��[�||@Lehä�'���. �?��&G�[�� �`=!]� �8��B�)�������D$��9�� ���������/_RS�D����@w�: ����*D":��t�@ʃ�	4���RG��~��r�D�"�
,泒rd2�c
�C �;��N�c��{HG�L��j�\w�� �r�cw։Fx^�����b�7;f�N�� ^�Uz�B���p�,�TV�-�g���t����䎴�{WB�<�;��~U*D�]��/�����������+,�CZh>u�Ћ��A�i���o
����Tlq��?���6m2J�pwX���x��)Y�d� (E�:8�%��ds���L�+��9�v:ɌC��\�k_�=; ����l�er���n� �ň;-���y*\xrz��s��0�KM��_�6�z�5u��:ro�m q�l�&�2��l&$��ϭMaf��rb�G���	/(gi���G����%K�߫���T}y<������"�-T�[J�R�wZ�i�/e�,C�����E��$Iٍ�J�dKb�%�����;��~�>����q?׼�y���|��9�C����� ���9���^;{���:��+�������K6Q��c<�*I7��8������)2��4SI�ϟ?�U^��a�3
ͦ(�����7��騕��ā}��-}}W���c�i �|�{��E:,� foG~6�K$��n�E
��)F�v<�T��%hB]x����^5Dw`A�L��ع�H4��K�>r65�C����ȥb$��1�V�j'����j6
[���.j����@߼�*QÎ�9�ub�;P2k��o�y���[n����Ҫ���P2"� �X��5o����))��=����z����ZAx�\�) ��T�%�W^\�vJ7x���^����C� ����K����8���*/\�ْ�m���'0ro�4]�����|�F����I��|��I^��ۚ�ߝ!� �r���n���})Q�f��>�_V-���w��������,�2�GYPr�_���5�!	|w P���|��^�]�¦IkV{~օ�����!���9�v�/��83��xn�O�Qh��Q��Q����|`U����9p�,e `�~�C7zW �ײ�"T�S �2���u(@<���M���Z���+��(�H�/402
����>4V�z�_6YtX�˳��\ 9,����k3PLc+�Y��7��L�SKi,�@r�����Z�~FF���>�i�*Ҝh"�����* �SG\A�㘟��O䞌�W��`_�k�oXpc���!�
G��������U���Gk˲�b*�sݵ���f��X��i ���f���R&Q�����|�?`�*<�Q�8Q�s{d�ζ��[�#�7zp:�lZ'������ߥ}��@j������_��}���պ��bY�e�K���3N�S�3z�r�k7�-٠KL)��%���>G���I�߸XPZ��%�����<�W��$�E���0��m���$����w.�����c�3���.�iL�gܡ����		HƏ�:�$R���_R�>j��И(���]��P���WW���22{�]�����k��?&���{{�}&�2�7a�7�C�o�y"�O�k�����ϙϢ�g���gu�31��������m9]��'�,�`q���	_��JZ/*2��?3uP{ye�t=n'� �8�&�̅�5t��Q[�p�b;tU��P�x��`���: �"�ܬ �[�n�
���~N4���|X�rp襤$�;�$8I��`K��J�ы����P�&	%	(x@��+����a��?�vV��E�*%���3L�����U�#Nhc���������d�+v;.�M�8x���l;RN��9gD���Kb0?�����cB�B���݂"}���y�˗�AvY��I�[`�E�KF3)۴��W��7�st[���+%-O��%���q���E@=�����.^��?���6  ���@?B��"ŧDJio��wsA�6� R��(�"�_V��� <f����Ԋ;-.,lk �ӵ����@�$D�����ؙysl��3���p��oq��>�3�;���g�#��Ř2?A���_�g`��B�h�q���ͫh#W�g���z���6�d?"N����ԭY/�P+)L?iZ@I��D�R�vت�N�hj��0��p��¶��̬�ο*��m�=�^����$�����?�K�6޳����TV������;4��-��.ԩRz�R�G�BA�;8@'���z�aˢ�I|d�A���{C n��ٱc��/,�~�zK]�us�B�V���b�L@&PY-���nu��3a�W ������|,�3���8���[�D%��/(,L��`Y�d$���b�
�Z�37��CU y��(M��X���B[��*ɘ/� n�"�޹sg7����*3�ALIkx�������N����~������k��l�3���M	S��"�V�c�V��� �`]΄^�ĭ�R&����`��{�8��+���_�Uͼ����|6�L8���*�|e����B�Xh!'/oG���n�.�O]��##�h�Q��G��Яԫ�Ge�����]2�ެ?%�o��8ۏ�N�q`ǩ�[r����������u;��ݏc��G	WM��؈�T�ȍ����%��p�X�D���䈎��ݙ:fw���	��y]�)�\��"X;d~]��V�Y ҧ��V㎮&n�A Aibbb�ڏE��9�ј��ב���Q��ޜ�s`Ν[��,�a��d� ���������s�c}_VN.�;������]t`d�����͵��<0d���,����۩;�Ilƈ2Ͽ��!���$c6�RQ���:\Y����i����=�W9Y~�'"){u�.HQ�Y���T�L�z\�X����r܁�$*��N��T*Fg����uq��B�;s���ukx-���{0�9�����H����� 1`V�w�"���c:�����sQ�Njg��=��Nk�)y>@D�ImmW��ֿ_��rA`�c���̏������ܬ�m�����R����T�jy�S2*��#��m�ɣ$h�l�w�DL�� � �|����ɴ�G�*l��cE�Vw��\[���6E����N�gY���vz,�_U\���LS���H�ވ��JR�
�5
�P"�e���R~�ֿ����8��*m||<���:�����$�E)��h��xwi���z�FA���ً��0� ���ZW��=�c�j�R00!�L�?��):�T���������'�0��D��9�x�L6�} O�d���?S+Ʋ$��h�ಙ:D���O����S4��t0�$B���(���x�B���_Kk�i��En@䥯��č�����6%���D"igt����ö���l �����>��|}����ZJ؃�`�e~旕�.�v>��>�8���n�_,BI�����y`fiW�_4?��,O�ymzz����:�s�Q_y+`h������j�e.�%���ϒD]a��U�Ev5�ѥ_/+��X�w#�q?�?��0� o�c�K���)C$Nu�����r�a��誯r��n�-<���Uz���澖�PC�T:uj;GRjj*Z-��	<ah��{���g<�;������_�VV����C����.�����e��Y��l����-s����T�n[aa�j�X�Я9dJ!e�>��Im#-VFa�+j��y2nv�#���ѣ�w[G;�dK�2�.uR������~�0�A8��#����nmpU��@=��2�$q|�$���O���Gդ��R��:ܡJ-e��'T���d4n�X)��Ϸd�W�����k:�n`c�w����g��J�;�����
"dj9��;�x��������t%w2� ����_��++J�DϠyE�2��T�0��
Jy���
ߓ�Ri�,p�w���XH�ιћ�=d���ٙfex����*��9\�])�P�f���M��+����������M����,5�rN��F�B���퓬����墢�Mӿ�c�ֺ��~6�{��/?)¬"�E�u2�~�����_)��F�����H��7����$�E���<8��P�2�KNYW�KiSo"�vo�o������}�Z<����##�k��P^�<#F����نJ�����Y�FP�����!�>w??1|���d�}���9��\,BS�:��LW�z�C�ω�=G ���簄�����R����+�|_{�=X�&?1���b
���Ĵ�����ʄM�}�,%1����܏1n�5��AW������s�t:��@�2���B j|!�{�~�_ɚqBYx%P۸vх�=�ɽ�S��z��"����lQF���<QY��T(D��G�P��N��'�$ŽE�%��@5������~0`�� +�<R�3VD=T?�(�2����&��i�Lu�������Ct���V�ж\@�����Q���� ��\u���e.�ڏ��!�x�E"�Qi�"��+Ɠk�:�
�	��ںA�'�j�!�}#�6�6)�%`yn�5RIz/0}X�LO�]�@1����J�.�&i}v*5R^���/%�fTc��6���6�]s�4؆�x��!�O���p�-���1=}Jݰ]������߂8��&8��xv��s�q�����˫�ʎ���5f���ҍ&������*!�6H
�c,l��^��m�1I?��#�ϟmH�?Pߔt�~�Ȥ�Wq?~���sR�j���44�w��42;Ǔ5Rl��֯�!��U��8L��d����ĩ {�{lIR��lnp���D}�)�f_��'��J���ބ���澒A���������%�$��tٙ)��:�yiq8)ȹ���]�и(�җ]���W�r�eHr<���KS��@A����ɘ������J���u]���d��$�>��l123ܬZ�U��:v�{�h^o���ࢎl8ux�A�.TEF�(Y���#'*9���l��(��t9J���4{xe@ye?������8r��[=)�l�R�屳�i�^y?^� 'x ��4�Q�y���7@�IJ�x{�3��5ўY8I�3]ڕ��.aߥ?C����~w�8-t�<��ԉ���kW���r��L�g�م����b/�5�_�,�g�[UA~�����;���Y��A�G� �"�..>>>٨�%�ڋ�)�=�!�(�ms��W�A޲���q_ ����`|Nr7Z�zB�;^us�2cE_������%�����P��d�ֽB��\JT�-z줏7��:m��1�83� ��p�/#�t��zb#�ՊJ��o���h�@�Qh����� �铼:���!/��9͔%�<��S��C��m��9�_	y$j�˘�U��%�q���^
 ��ڀ��1�w��t��N�V����`c�\051auj?�I`�$�ךD����]��N#'��<��-�� ��,�{����:?�[�wnA#CE�P�����ٝ'4�>�XV����0�X>{����|[�v�1{���z���8^��,���7��ח�ߗ��&k����:�-�p.�&�/+�u6�򬋴 �����\���Fя�r�3���u�^����w_^�)�� ;6�]�یc/Ľa��?)3��I�Iz�A�h���N���F8�e'���r�˜+]z��D@#�I{���`�Ol�Ь�R�8;U铣�)�K0�c���8!�3�N�{�'i{9̌���o!eft��Du�J�|o��N�"0`d�/��A�vv?��{ovb����uoH��ot�CV������\�EuǛ�e����Z��Bu b^B�����AbVS�ZTo�x�ڲ���*��o������ �%�$(㿢���xHT)���p`c�kk%������1>""�=�1�R�$��������?��і@T ލ]����b1B.uW�8��8����W�8�c�-�T���J���^�BlkaVJf�|�m�R�����ij/��T����2d��W�N<�%�	[�׃)~����fff����Yp*Hӑ��$�C�XȞ���_]����Bޓ!��x�:/"�FU�ߖ�MMk�@u�OZ0����c���cJ�8uXc� --��9�m �
�*r������Xwӻ�P��� �T��L9l���@)��$��(��3��� ��r;���6��>�VD@�W8����}=���}N+�G'���V����UTD����!�!E�C���B���7�֊ew�[NO8�G�f�ᴑ��q�|]��hD\Ee ��f�<�?�ro �ڐ��%Qc��6W����)A@�N��Rau+5��X߂��*Լ�4!�����6��s.9���l�H�f^�ơ=�X���]��nҐS@��k�ϼ�8�Xd��$�!��Z�~����<�1�	��pQq���J"��F<��=��XQ�Qhr�=�Źxg�H��:Lلi�~<�^���=��/X��n}�dI̡z`(9ȎVӧ\��)� SX����`E��2`�?-.\Ml��VJ��#�<i7.��}�|6���X�~I�1���s����`;�b�u2ɾ�J#�����%��R�J�K���?m�i��l(����3Z�WQI�x�����TG��7&CscM�i��!���*�7C�]Z%��n=��v�}��;����N�@D��t�&LB�Y�
�
L��y����4�gј��q%�����ܖOxmy��5�����O~�;~<p.Ր~��������ST��˪��e��[���.�ۍ�I��<��Gm�4ʓ��;��FΔ�X1�wt�ب��YxAM�2�bI�խ�c��#1��G7�i%�u�M�E�6�ٙ���A�S�I3Ӧ��X'��������)D��YΦ��\�s7,XL^�����������BuA�9Ρ����~h���I���_WlHR@���Ȱ5�<�<��ʽ��d����&a���r{��h�4&O|��1qarb��R=p�*�Ἓ�(&o��a��l��j��e�/����'���H�?��Wo�M�#/,�<�6���,�1y`���-��O u���� ���a�><�fZ\���RohIY Um�"�q(do0�t�S��^�ܜ�1��� m`�и�5 ���cT8���x?c���}!	ǜ0]k� R��X܏�d�c2���Ol��&"��qr�L�$/�ct��6ϓ\��h��S��]��X�`t�)��:L�>�M���l�:48{p�w\P���4\���D�(���?�|Ĥ�Fhbq_������X��_���V���5^0=����"��O�\�hI2Y��P6G0/�*PXd��K�z��Q�	?w��II�]�/�]� �'k����0��^�0��+j��P%�;�B��j+�f۬��*��a�����z6U��E�w���"\�v���j0cf�Uݠ���R��@��U`ldٶ ���b�����b�2@2Т�X��l���*��OYI����<k��Y�6����L��l�P}o:��u	�	��ͰX_�.�SމΑf:�쳶��~Oҙa�<Y�9XZ�����L��&�<4�Ί�[��|�e�G�k��?$��~������z��um�!�Q���T��@�=IW�<b�[��� y%n/�,m�<�eo�&4�H���@TN��_����k�С�V6��`�_h`�S��&�o���.{�|�3	G���К�fh}8�~�]/�A����p� ^���u:���xZ.��Q�z��A�¶�(s	���2[0�=+��ht6��#�8��l��C�3A{%$��;���'�� P ,��s�=�4����?�RL�$��N&� �SZy&f sF�e�.������,�VO`p�
��r�BrĄ�p
?L�D�d���e���=�U�kD9o�}s�X����"r�}T�*�8S��>�Q���;�E����76�A��,�ʓ�6���o1o���Y���)AY٦�>��՘ͱ��$�cCBYו�zG���S��İG��&`��`<� �O�L�"!�6^[SV�&ÕȓA�o���bʻ�!O��!��)�'��m�O�11Hm+���d���4�lR%�������'��DQ6L>�~#uy�=ɫ`����m�H���"����
�6�4�@%�_��ʌ)+��<s^�&l@��=�fbzÇm1g�rڀi�o�T� FCm��l\wz�"�V~�#p��nd���L�Q��x��O�q���_[���8��i��Y蹻��3y�����=�XlH�4{�R�B�'��&J{T�6�JT�.:H�^$*�u*���.N��<��0B�Oڏ���~y�Ӂr�:`mY�ɢ����itn�)c�W�*a�/�M�_�9�4��5"sF��x�)�݃�,��@,�A����0 S���m��o)lb:u�;;��T!�qe�:P��0�R�nܩ��!!)OI _ܸ��I���[�AL��Zv�xx�G���Ïd٬�SЫv��{m�����Q[5����;�3Ά��$�U	<E�X]H=��1�7�ڞ��8��j�Y�٠5���|q�`-�A�������I���K��0����q��[	��8m�!,`�x�o�;3}4^�
:��ޞ��'��V��ul-��D岀�ڝ�C��'C��>$f���ěP����<��'�t�e/����:���D���*���BY���ݫ�IL���y��;�l&�2�,�m���M��z��VIܽR���(o�p�WR�^�� �&�� t�� / � �Oӗ��|6C�C��;7�\B�^�#@���f{|�Z���G�V���E��SL_	{Vvψ�)s�Pr(���(8�v+�W�#��G�!��q�֠��zІzw b�t���N2�v��{c���� ^�z����)�'o��U���[���F}[`eCZ�V4�7߂���N=�X��'�v�U9�����eFu��13�P
 諥h3E��Q��}?��^�/�h�G�όTfO��Jr	�

8)�ߵ̫{$���\���:]OT?Y��W7qY���4�K i����{�x@p��Sf���O��0Y6H�.$m�Ѳ��gY�-��t��v7�7��m8��\� ;����C��J�[%q��
����@EH��,�YEc��|��������ʯ�"P nbbB����YT�c�*�M�T;��������T��Z�#���s���'��nGc2�X��ee~�z����Q��3k)�%wv�ƞi����3u)h��缄��a �cH���U�|~����+�B;n�ً�������6�"3��ȌUR�BS<�nX�o"� ��٭t��l~��1�������k��w�f�y����5� HK�� SOI���2���ܘN�S��y��xex�M��(�f��.��
v�D��U�ۻ�����y�5N��b��LU?�����G��B��t��C_s2qݦ�N9X�Hy 2����}=��B�nwO���xR3�2�#�������w�ѷ��x�vU	��nn�k�x���(��4n��m��Lh��e����o6�`�"��t���Z�m�a�
��ǹq �E�GQ��7w�cu�Ȳk��̻J�+�n�(���<�z���0�@�H1�G��z,H&�K�گP����?B�SGg���&+.]Q_��/���0a��t��� )mC����˙�f�б8ߜ�=;�M�hGp?*�=#܇6�(������u2yҼ}�Z���7�6kE3�:�w�����y������&��II?���,*�BR�-S�L��/kr�x�=��=�Ӈ7���7���!�N "�5Y��
���q�cQ�bz.�����pu�@*�3?���B�W�P�hAΫ$ړ(sFFF�u�͋�7K�~#?k�����s�ʼ�}����MB>�um.g�Q�@ٲ�hx4'�:�Ƭ�uV2r�d�n�X��=��Dc|��
��;J���Gާ95�*��J3d��,�lk��,̲r������/���T'���<�m�v����eh�P6�S��,5^�s���hy�"T�7#1��JW�E��jWn���Es���7�ˤ�gF�9T�h���S��̏�n��*zif���С�����E	tX�����q�����ĭӿ�t�,�19Q49��XF��'� ����4V�dsf$T�a���� �q�3�D��Σ7�&k�(n�!l5��\�ST{p(=�XH�I:���ӯ@E	]��f|%Q�m]�����4eש�i�������8-�啊VNf��:s;���"�C�d���U����kʵ5�B�Q]�!�-���+�wb����g���8��[�� �C2�xz��y�֍���-=�m�u�l3폳�Q2%C.+w���z�M�7�@��,N=���=)���&lW�!��H��(����K�Bu'���g���O�;�G�G�ib��ӧp���~��ӿ{0(J�8���sGG����/���ˍl4H����.�ߏ��Ө��&1�h���������5 r���H��+�)���A����ݯ���ո��L�s�	���\b}��z�P5�cD�ݶ!3����<�N��n)[]�"��������ow��V������?fİ��3���X�o_��No,�}�8�8�|�Q���9Oϸ|%ݣ@6Ѿ ��GI��{jb�]?�G�p�UD����u�M.�9��%_�� αj�S��z���t>lX������&��tvf�����cO��͑8��.�q������){�b��ᑏ�����Dr�[��$E����0;�CJZ�:���YE��͋�>�)�6#F�b��Y+ �{Bpg�p�'�M_��w߿@�T������77��oZ�����0���hYl�5�5�]��yUB�]'��{�/^��$Ts�kE��񪌴�'�����Y�Y{��°_��:(����k�Y��b~���Đj�*gE��!^�>�Kp���j.�6�*$,��!#�f�|����3{ �9W�R�b㐾�{Y��^�xŁR�7'��W1,Ck��d˩ix&xC+�W��h��C�����d�q�&�.� ���͈��	�������)�U��e;��G�7;�E<#n9��2�����(��B�~&)�q����56�	���*�|����c��fҧ�zi����'C3���"�4���H�A�$΁'��$����s^�\���q��@��]���^����t8U�~^tA�W^���������:$��������\ڲX_3���V9[N
��EB����~�-�B��b�h����osLK9���x�dj��4o��&��)������}���D/����������6�M�^x-aL�,R�p.�2셈��km'�����뱏{����Xa�e�`�k	ҙ������ShE����~[�`��p�p�>v��
n��Avû�n�u��T"z�^�����4Ϻ ��Zj�j�3�]�Y`�#�~�k�6'$�M���heu�A��JV9�H�j`w����caV����n�P��
�t��P�N�����r}��@�� Cq�q�š��q15jU����g�����z�I��v����Qi��q?8 ���#��f�r�Z�&d�jJ������������;4"�-��a���S���u�}_�h���߬�𣀒x>�(��wr�eM�-=�c2�ǰ|uP#��1���^ci�p׺91,M+������񰷒�O*\A�.(��`�E�S9�^qq1�� �a�gb�.�r��CW�u���t�(��"E��P|���NHI�>��L2��۔;ZL���N6��&�,��3g��#M�g�[[[=��a'�sv�����x�.���ܬr�:44�l��͹CE�j�b��Ĥ�7|�v��"��v8����^l�g�S���.�d4�, @"�#�>u����O���ZE;i�L���ߨ#���ɟ����0���p��r �YBBl�X�����:fy��0V������cMk�׃��$�t�a#�2r���#o��z���Pxn��BUH^S�L1C5����R,�s�r)///;X��-t��O�0~��m{��	�Y4��ۤ3A<�]��~��5��U�P�������h�α��okD�ɡwT������ѡ��0!�Zԛ��JօG��9���&&F1�|���^TQ���4��t6v{��o����?r�C��X�j��S;VZ���2%����]K�w�7ڔ;��(c�-d�`���hoon���eq&W%��G՜!W�E�ٔ�����M�E�rhx��g����T$5�.�Nj��ѫ�L�=����u9"V��,=�tPIF��t���Ӡ$���Hd\2����p(�F�M�X<S��w���[��/;;��]NWk���b�]�>;������GX�K#��f�c��55�?jQ{�������������u��U�����K���/`�e�b�Jx�c�F��kڪ����D?�ځ��Y�Tq�U���ǋ�n�]B�H�H�2[���Y���ү������8h����R/��v�֪���$r�^�4;�`�Y>rW����o�Ӂ��1�8栏����<���4�$����|���u��?�oV�}�����>��M�.4�N����� xr~@pu7X�@Q�[����(� �d�q@�\L�ʱu+�&Q������P���+���W:������<3�ް�q������)�=M�»��U.��:&���_���ϻ�A(&s�v.���A�&��D"'��?{�����0�eR`�u6F�\23��+!��_������on�|�c��T�m�=�d���f^`	�5<<�K$�.�b�]p��{�>k�s��+??�v��¼�r�ҥK�n��iVy��*t2{���~Z�zy�AwWɸ���x����
��S�h��6)���iL��Q�ʤ��}���kv���F���傂��٣�!"K��������I҃Dy�S�MP{1���Z�b���Cvl����7��� ;7��������_���8�*��m�:I�ww�8�S�������P�q㒝�s{�o����L7��=��0���"oU1n߿_�O)0�6�\۱cGpm%p�E8��C����_���{f.j��9`.?����'�CBd9���㵄���bss���i�a'~x�Y�ۯ/{@�q��jzj�ڋ��.�^�Hܨ�Al� [�����ϸ��mb�H�BK�,wJ	�v���7������v�W��Q���+��2�V�鼶?y'Ļ4�
����o��R!ȩ�������o���ճ-�m
�ܞZY���b�3u�-�R7���",�r�WP0"!!A�e��*�jz�X+�G2�W��Ш��J�#�=��8d���}����=�8����חObi�� �����D�FF���I������yфx����z>��'*�2�"��+;��9���	>.$�:�Y�;�!�t��;������.e�^�?�22��2��9���!yW�p�h;�p�0&n����m�^�q��oK��2͇f9��e�Ёq�ʻ��b�l:}�����f>�t��qo<)-���H�y���t�'�V�H��u�!<b��z���`t�QV�m�c���q���5yN3A�e�ZM8ܧ�~��[��.$�ʹNS�ed�F��>�t#�@C����5qN[���7??�rq��uL��)�l^ǣ6S_4V�SUt��i6<-X�w���%��4;I�۱�ʛ�c���⭭h��E�k4[W���h}�ֿ`9bp92.?���4kiR�Z�#�`fY*�;!W�#�ZQ'y}��"`���1�Kre*Xy�hG}
}�M�A,�I\�Җ��ぇ+�jii��ż��bM���ZFǖ���昃�R�zNSH�6�ʎJ=_12�P����3�_���ط�]]��G�4�0������A�Q�U����YO/WT䇷⵾��r�#�lM��${*f*�aÆC#"�wG�R��}�ά8�#7�@���&d��Æ���j�QWa3�mHI��w�_+++�13�@c*���.�Y�X%Dj&(y�9N�	]�ٍ��KO�U� im�U�yx�<*O�VLz��su����l���\����JɏM+�bM݁�e��Y�;�Ka����T�X�p�V��Gbbc�\� �}[Bn~\�ԃU.[�66�:�Iml�}q�*%Ѭ�wiJ�����+�h�R1�>�����2�\V��$����p.���I�v���G� zwg$��!��U����ܗ/�]}���^z�,.+���)��8���Hv�C!�����I���{Æ�I3#_��]j5�pe� 0唗�֒�4K�c��/���M�0�
{{��{��z������`S,mE��h�#+[�t���.UN����K�M���T"o�q���������]r����������]\1��J�tL: r���ݙ:���yY�Zϔ�=yyޠ�d�3����_^{|���KD@�T*U�'���z�e��^��9��F������ҥ���㕦H��T�cJ�& .ɞ�V�]��B�Mf�ʹ��䍍ud �j���o{c��x�`0�W`������j%�&:>M�=_�Oa�~��G��鰪3�y/ ���H�h�M��d�W�����a���ҳ��qhO��9�H1���,�wH0[�s�rD����JF�g�t#�e�V��+��=}�݃&�qZ坦/_6�\{k�ܠy`�Ɋ#��� �n��w�q%�)�B�):�=�{�����
��T��)��]�n��XF��Uҕ4N��<~@lK3�� �7�]��:���!,� ~�!ϛ�j��Ex��XN�������XUG(����N�zF��q��4�`����4��3��]���������8��H����^^r���Kۋ:m��W�:�����'�s0J=ʉ��J>����E��m��ۿ���\�$�&<ss�ZV�y��KEn�ׅ��`��/sY��x�@a��㲋쁌��X���Q��ײ��`#�S�ԩ��#�AD�R�d����U�\���̳���?�����_O��q�$D��3�@�&H�Q�����ga[J| !�7�}�i�"�.�h7?�E ��K7�v�A��W�L5s<�������3%��F��3��� I�(��taG��m�M����M�%��fܢ:b��������'�ee�͑2�%�}�Ŗ�X��c �W�#�F΁��5��֦J"��i&k�ۋ�� ;j��Ｏ��G��{�#m\�J����1���N�.�jT%1I�я8�	{�!��
��ݒ ~�,�X�0�W*Ôo4-ў��������I�G��"R{
��Z�^(��g
7�A29��if�C��5�/6Y�K���AY��#Қ0� [mff�?++�+���z\����n��a(2��tD��]��w�DA&~M�!)��h��N�{�����#���|�������y>�_�����-�>O�@�SY|�r{S�[���zGЫke!�BRG:F����GMJ�N���������ٟ'Zoom���Ze��=�?{ձR�����T��W5~M�J4u	i�R'n���&
�KK1Zw���st)���qܤl���/8{�,J;/��^;nP���X�0����'7�Ď�܂��a���d|:/�e�ŷ��g I~5k0?���|�+ �.���/ij8\�����)�~FG`��Q���֑��忔�'|,��l		x���H�,;�`��g��'�(�%{V���n��v,Rz5L6��|c{����J^ l"!��,���.JSw���0f(����H䐸zt{տ𷅹��L��җ/_R��F��pN�G�-��J;|N����
��K�=z��S
�\���%=�TJII u�g����x��6�ia8#kj��á6��\���&�� ���_�==F=~�#D�s~��>�e�6*�x#���x
����D ��E�Q��>϶��G�屙r���z �����oL���Er�����mv���0�B�^�|��E�NQ��)9`��gvnaa��R��;��l�O�>M�GI>3�H�jP����jN7 ���6?q�g%�  ��!o,���	��F[�<s�}	����e(�m+��@��c���}�a�"~�c�$�S��.�'v?��D��Æia�(�E�#�(�� �/6��:����״ �{��W^W"Z_V���(����)��/~����� 6E��ّ����a �Z-�p}o/��Ԍ������~-��~�n�j�BؖC9)\�<��?�pȀ��g��{����1Nz�S�P�'�*��b����~tJQ���Cf��L�m�9�]V�i| ؆r���(��&4��ʈ�/\5������Y�w(I��=���5\/���݌�ia�,{�D..6�b�U�"�`יe��(M�y�)��bp7��OQ�.�SU�-�N;�.�ƈ2 ���χ�	d�&�)�8�-L-E�b�n�O�ʡ5�A��y��p7��������2���9�ŋ� �%F�>*�pRW�����|-�'�ˎ���%����{�踆�%q83$���@)/,���[��
�*_��+�^���2OqH5ҟ��O>���"��{�DX��O������h�TS�x�ï^�6�����Z��}o޼1��Oprr���RnY��j�{�*&�F��^�}[��!~Jy�Z���M
>�4��~]�0t�1�捝M�KU��w��h����0^ �ZD�?�'���w�똽�m�]�^Q}O�1�2Cw��b�pz�L��-X�|���D<���Y�	q/��T�N9g�M4_+aO����C;�RݑYo�qps�C�%��!50^"Ja4���uX�%F���O���N!*��x�<J�y=��z�y@OW��Z|!v�auu5q���+�4:���C����ϣ����b��X���;�hzO��Y�WD����~������7��t�wE	v\��14���
Ѭi�	�V\�ʇ��@.b��|���0��B�h�m~��V�΂~?���+͸�|��1��AF����jhd�$��g�3�;�2� r�D��C���jG{a�]R�2��C�=������WrwX'��~�ʆ BD����q����y|����I�;;,4�ӏz?���ka�������m�W��������]�&��%E��dP{����B�|�	���.���y�&��a�+���E%�L65a��g�S�b��z�w���\��BS��� �����6F��-i��?���AE�v�}��f���O潀@�Q�m�bj�xE�)�Ӽ��fD�C�n��c�σ(X��^��N괺� �uѫ�(�G�T��K�AO��2n,����)UF^}xƥ��B�=����)���S	�"���0+ .��6�VUU=C���y����7y)&iE�l�y�\U���z�,���A��vE ��\Jǣ�\��IqqȦ6d��@���0���� ^����2���y��Wj�L���u\��[�����Wr��ݿU ���jI��3Vv�-c\K;��t�e�/<lM)���4 _)7�_rq��G�%��g�(�13`;���y�C�g? ��Q$XYY�w�Y��h��F�\�Y�b:1D�C	�o��j�A6M�'i�ޝ�Vg����	���4�c��V��=R<C�ڗu+�����;� �"w\j���wG��ёr ��m�=lq��!�F^�ґ��UJ�^<�5ڞƵ|6�:D�X>��y���Uz���_�͝�I�M���!��IF~�={���-��4䅎G {m�!����������W�vj�a�z�;�?�&u�+�`PS�l䧢#\��jD����E���P-��loXx�Z��˗�}鸵�����~�E�# �y����?���e�'!r���_�7G��]M��S�������� \| ?�x��������P�&ž���Y�5ν����z{H4���-��D|Sri�~u��I�~���{<����z��OtU�/�����<�".�!��'?U��CU�͌�����г����q�P;#m�s�����x�ϡ 1nG�蠒
��8����]����E�Ͷ�ҡ��R+���9U��j�4�V߁T�����w������Gg����-0{yz��cw�w3�R>�x) qvo C��6�zj�E�i�{��t�� ���wmफ़6���"v�bz�A�0��1]kuVk=]@�.�A�������XA�p�m��rG�P;�/E����P�KllFOdu���?E $:��쭵��z���n�oca`�*V�N�"�!���r>1]��V.���x-�e��3�<�gb�e�Q7��	,�y�F�{�g0$u=]«�`O��X�I��d�&D{�AJa7n���z��S��A֞L ��CgK��6ݿoZ��5}��m��,�SŞ���SFX'����rr:)���Ew{��������s{��|�)��/s0S�[u��\����}ny�2��;&�����p��繒J}к�Hf0T$��$��M)�#�g��)�C�ft$��NE����ds�8F*���#��u�i���g_�1����K�)/K�%�h���D��嗊��R��ɑ��%uJ�e����:����q�wG�B�Q7ڻ@�2�:�|��EIBb���`�#R��������s
y\��C�����XVq����fj��RUcj`-1����BF�#��M5:M��b����KГsG�	#YlGy�Zn���?c�3U��$�m��a���XF�+�N*(xɴ���+��ŶF�2Y���P��h!��Y��D^^ސ�4����uZ/������uR�^X�ӏ̞̓hO�۟e�5��}�,Ak6t���`�E:Z���g����p9��v	#���J.\0�$��;퍑��..ೡ{`0���UA��A�q1�M\������VD��5��H���J@�āv���#f<W�,z�O���>��U���^I�̅�i�}��򽰹�aA��u8���zX�����H�E�j�Y���/J���X�o�����{��}Tva�<�gH��n�{?8�*%?��$^�P�+��BCw�[�\��mQ��D<%%��)���j��|;���ȏ�ߨ�+�dD`���=Ez�i ���"I���k�I�䙨4566�����}�a�%�|�Y�D/!�(�?�]�Um����Nq�P�0�_��Ե4�͡���J�)��?�v�����4�K�Q��1(�^��wl'�AB�_B�M���T���V�-�L���Zڏ���p!��d��������y��^�i�7�������շ�T��%W�Wفߋ�gZ[�oj^> $U�0��j ᷴ\�D Z� rAqq�2>��fyYA>���1����2��z�>u�Q,=9z�%�����)J���b%�e��)⳿q���춶	>\ՠR�0/W�i��e"��	�p/�B����zϸ&��ׂ�ւ� �*"E��ܵ�a�H����k(�
����&�P�Ћ�KH�H�Pߙ;���߻�8�}�s]י33}k�V�ܹc��'�C&D���^�tt�>RFqQQQK (��<p�1d)��Waq��N��Ӄ��%3yc�����[q
0&���]�6$�B�+���D�'�Zk�K9���$c�'/���4S|�K[����:oC�}���U+ ?�K� *�,����¬I L�_�o7��5Z���6����b��_�XS�k����~?lyF��zlV��^sɹ�)�[4n���Z��k��~zO��-�h�1��PP�k��p�nw��-�F6GG���m_g���H3�~>�wlG2��w\ұ�8�Ky���'GGG�����h�������Z���|���)z�W��J�oSuc>2ʠR�����k���e���^02��^�0�z&�9�@�o̩�,�7݂is��g�P��< �F��ej�ǐW�_�%���JϺ��8�7��B�HAs'ô\gm@�٫K1���ȓ����[}.���=(+�U FŪ!."�9�r��)���9�	��Z��ص����D��������?J���c�q��)��Z�����F.�g՘���8]�j�c�JIL|�|����������?mA�Ţ)�?��V���������! M9��d=�A�6��)��_q���y�k��F��öf�+m<t(�]�5��	Tv0�@�]q�Q��b�/���vt� h�Ĥ���v�m�(?o��(����ʍ��,���wA��	�|G9:�֓
��n�=��ܡ4���<�c����A���8 �$��h���ic���Hn�u[����g,�`C��s�۷�[{�Š$����c1A�L���N�
������2����GNN�`z��ii.tk����B�W�W�\,yWR|
6Uмe�e�v��h�-O��S�ƬTBT?�������:�������8c'*�ɩrX��8K��C)q���$!�@��T��B���U����*Ӛ*�
��ogu�LY>}��;u����=�Z�U�Q�M�[�f8��G+2���7������A+~�����n�0�+)I�@y%8��[�\���kH����:�K������N���1a��0zӬ�P��_�\_�wW"�Dq�G/}���i�
�7\��O�r�{8�d��7K�.���%V�
>�٢�v���+���ަ�������e֤h.Fɩ�A��Ɩm2XWd�o���S}�����(�²�nd�U�\�o_�#'$$DJ�)��nhY���EP�~V��fL�x\XD����w���� �#SK�}d�a��'ON.�%��Q�$���A�0��)��(Q���6<�đ���i@x)ӭ��ܢ�i��ɯDxD��ç��@q��NHR$r?"(�.�^
m������P�糪�lD����B����nR|����e����3&T��X+����*�9w�K��k�n�,�@��dpYF�JA����"|/+'*N)�g$��0�hR�w[c�m�ې�Q�έH9]����o�1�ӯ�m�J�X__�y6i=���D��+�:5��������*cmm��ί�/W���Q��(� ꙄĶ�v��['�	������!��P�m�<��c5\����p%y���W��w!k�Y��v||������2<&��hU��B6�������YO�&ŕX�D�#�w:M�y�"7�����<z���"���EŲ=�����]n\����IFf���;�|�maF(2�+iq�6ſt;�;�]['%�	�B�iZ�VJ�l�n��m�0p���ϻ��9��p0a$>��N�%��۔���l	
�����.
f�+a��Uޞ%uuJB*G��MM$`��D��H�s�����[ޭ/�[Α�1�_�|�G�ZD(����BZ�3���J�v��0�\`�>��f�2{i1\��|�3A
�D yHFknn�@h����e<x�@���b��'��LMH H�Q煈I燵u����Ng�꟎�\ˢb��1���3���c�P��(��荑�	�+�<������=����>�0bî�$�UJ3����!�E��Ld��[��nʎ����A�|\[�ͫ��N��x��X�uII@B���7���y�ù~U-0x���b겻�u�,oA��?� �;��}��c���� (���&�0U����"�fOkt���}��z�����Ik~��@kk��LGGW0#'xm=<<������/dׯw(4�<��E�`A������j��2�����c��J_q!5�}d y@x�SCl1�d/+5�l�P�����ׯ?h����V����E"��>0ʑ�V���b�P{ �b��i>PPPp�v=���"}h�o $v��V��r"f,�:2v��r��Ç!rO�G��Ua�!~$ߤ�
�~p� �XUU��������=�
�̜�΋.6��ͧ���vvv�~4��oC�}�H�4���˗?���?���:�Ɩ���d����-c�.�Bj��Sx}L�Y���ZH�m�u�~l�O�E����<��ѡ��㺎��9Bi��s�?[�6��g�h�no�HCE��U6՜���N�`W�����0�eĽTYI��
I��'�m�g|4۸+@Dv����(�	.�]�2'�JN,�Y+E���%�$��:7g0q�,���!��% -?�BC���`&�p������-���8�J>=02TtI�z�+
�<@Vc�{���S�?�7}�TUU�8@�A��M}Y���=ո-#����Tɛ��ڪS<��f���m�����g�3�;���l���L�,.d��=F4t1;���԰Jz���#�cs���fL;Q&��b:C�(A�~��0V%��ff�C��e�����RGc���)}�cKGF�?(^R��ˑ���$�)]w����1��@ź����=�!�oB�T-�+��G:�K�u%�hю��3�l�ڳ���|�A�����O(//�ҍt��.���WE����r���Tav9#Í>S(�c{ן�� �!'0%�.i�6�V,?��>K�Be��tٵf���b1��Hk�6N�&����Y-� �쐪ͼ�Z�6�1E��t3������aa量&񴜰���jHQG��*,u��1��}�8�4뵕F�̢"���Gޜ_�;�k�͇���X��7�e�&�B�/ą�E��X�xJ
�/"�$�P�À*��2�l�o_����h�fĳ���E��Xe��h�3`Ŏ����T��4~-�!EVVVK,c�i&+`�V��3N��|�(�#&�4���9���3lmVq�;5���]Bq�$\NA���6;b�?�R3�;'�|>�~�@�]�o��F��X��ysO�I�sy���q8��f�R�j����%��1ԑ��v��Zi�t��2��-��Cq�$O�f�(*8Ɣ>)���#�J�[_zB�RAw�9�i��Vʮ�P^YY��C�������4��������g��
�q�Un޼���>,鄇� ��#ٺ9=��ќRN��k�cd�cW���89mmmfM�OBB!Zɸ����M���&��5S4�E��;�����gxx4�:����1�l~%]�RN�̩�ӗ��}��%YB@<�����@^���n�:W�A�Q��kmt��)4�|�-w�A�쬼�$�����͒=,�4�u#u��;�]Q�$��������˞����v0f^䍓u�q�Ȱ���o�o�xp4ŏ\	>��8s�O�{�=�߿?28�ۃ>V��������H�Y�d4��y�zy\�' Ȩ�.VL �Uza:+��'"�$�����rJJ�gr��3O z鈘)^�6EKl5��Ɖ� 	AyH&`9c飯��C�~�po���op0"&��j�y�dQ���A���%װ��W��ड़�o���E�ݬ����nA��$�bƏ���9��VvY\B<Z�{��}���5�(0!�"NǕ���(.HV���b�<�oIJ�A+� ڶ�&��P�+����}�Ws���D�U{���6M�9r�MU�ĉ�	"]�$�DN��ψ�ҏ^���	��W[�Ԝ��O�$��|���"�@Z1�V���c�_��~[|&%�-�-n?��l�qTTM��;/���h����LG*�6��	t�I��L��⯪i�(Bfx�j2εPu��wl���]�~u�W����-� ��<~� *� T! }�Z��>�Y�<�+66���Y���ZzD�j#1e�M5��իW���ˬ~	D��r��悁"	�B�u��<���l[p2s[g�۫'g�B'���o{����ށ�1�HҌ��q�3d�%�|������c�e>�o�� 7���53����C�z$�AKƘ� ��H}
lU�N�o�
���%�ups���d̖yc2�K�Ҕv���'�y�����:���,,��+��r���"/�x��Ux� ܬ��+�5lkJ��քkU2�R�o����[\T�5,�!������� ���"]�"����]��}�����<�d�.������>��ǟ���q��*S�S���*D"�a{�ak��MP��c�2�s'otcu	�_YSsr�{GG��R���>e�ֺ=�K�S_)H@�7����]�%��5������77�n�}����h�\���=�Õ:�
��?}�;x�˭=,���ȷ`��N�U� �@����OW��{���~H�`Ų�	 �aW���8�☤$uC��u-�������-�}��g~~^e����r$�c���[X(������Zdd���>w��DY��f@Jb�5�W� ����޵�V��ҡmiiY�8���7�����L�K6����&~F�W�2��-��iǸ`�B�'��
Y��F�KH���)O�L��c��+�=H���@\�J
%k��t��+�j����9� �Н���]*�h��Qᅛ��)�e��ռ�������b*c�#����ۆv)rrT1?MBCL���N��~�m*}[�X�?�X��J�crLM�A����ys_����1d�_X�f �/���`�c�����q�|��E��[Ю�h���"��J׶�R��XS �@mj]�Y�����օűj)A��VRIII�l�C{o6��9:;�"��#ZH��o���IM�Ԗ�a��U$/ݾf�>����MN��Z{��Su��wÂ۴��}�/織�A����k���}r��>��<�si$�拣���b�=eOҼ�,� �o��dJ)���a;��B�N"wl�&���8}�賰U��f�;�ǎ�����Z��ֽ��K?����uއ>+��5�~��k���K��g��<�iu��p덬��)o���X^$(Ү#�h�d��P���!�o@������
���5�O'�`kUi׭Bjii	���C��䦕G��v��D��#W�t�L�ԉ�>��B �� q����	�@	����A�d� �l�B�K�RĚgf:3�ۤ��J5�>����k�㦧����c��H��>�a1��D#Ci����۠��/.����[�	�$V������H/q;��KT\�+(Nux`��4
�9�.s�>n��"ww�iX���<O�I��&V��
�:�V"�(8X�d����PD|||��z1@s>'��I��j�����f�?mc�r�}�������c�U��*F�L���oJR���$ ��8�����f�6����p��Ȉ�מk1v��s��DE��_�J�:��O��=� �}r.3%��X!���_�l�"��v �8A=��\�a�zp��&�"}噶����#i���°���BΥ2�J-��(/�����A!9555{�]�����@r���~��y��r�I����C����!<�a��%v(��6~w�nG?�BĔ��722�s��U�t�3�;��5�5F��ż�?ڞ���Щ{x�e3��4�H%�jnu���Cc��8��驧;n*=x��O��Qy�2��K�5oA����e����=���^�{�t�J�l��P3H��̬���8�n~w�~r�ƺ<�j�Yx��}��'c��
���f���G��H����l�̱�Ȳ��${g��
'���{}�)/�����tM����KKK��q��Eᜐ�%���F�bP��@�����������K�5�쑏��ܝ]��_��b��07��?���ŖE��2��A�^� W턯���K r+%��z��vu�j΀���Ї������*��\������.&�^� w C{b���RN<��p1.��s Yw� �ĥ[ֆ("$���o�#DA���<�ٟHDev�S���[��?r�9!�j��h���V���t^XH ��c��A��Lz�u��T,�=t	�v[w��>��5���+7���ʯ�&1�����3���m��66�$�=���e&RD�̸��3O���c�nw�P��c�{e�9[���=��S�Q��=���N�s���B���r�u!�*���U�u�YXvw���S���P(0���8�8~��Qg4���Z����{�$	hV�Z�;E�(�-_.჊��}�jg%�V}�] �.�Ω�b�1�/���wGK/��2K䱾j��̒? �R4-�t��`�Ѳ�P�C������� �^P "t�h�4��D�JW�7��R�0���m�j���<��맮n��}���d/+������a:�NLA�ܩ|`���(�1����l���v=��6�6��V)�]��5�S������ξ�5���dO�ʬؗ5P�oc#Y'�"�����z�18�����^��i��.đ�2��L<�U�T��S� Wn���Wd�8��ӭ��~�(���4���ʝ��w��y�9��Ǽ=L�8V�_����ܹs����N)r�Ez�K���Jc�4 V k�5��R��M�C��.��� jf�4ab�����F[�v��6�������#@��=�������b�����]M�"Q�h�������9���:��@/��(X�ia��j�ȟ���MV��n�d)��rOOː7��?K���Mz�����GMϴ^�\��̈b_X�����!��ժ1��a��#��>���*�;�����Oyb��)S0"���ו��&���R��9�����9��]�$ Y��?fP�$�]]�P]�+'#7�F���תO�\W� �C���K�9��B��h����{�S2 �p^�A0W�NT0O&`�۠����0|Z��닕������RHI#1I>�un�90�A�@LnF�e�-���f�r#`��s���`�"r�f�	�5��\W�D��C���.կWJ' ��4=*Ϩ\�~ �pg�ޏ�=9yy�;ۛ�;��/�/�Ϸ¢[P�bNѾz��g���A��:.�,�������0��9�
�����f����R1(��=�O��ne�nRi&���=ֱ��e�ak�y�PՆ�$�<�u�~�FI�پ�\���/)r�hRQV��Z]�!�`X�,SZF�j�G�HĤ}���1����7���G,��@�����͸��!5,;-�fH|��dם]�� ����v��O�v���k]_&��� n��f��Ҧ!p���'��V�6��<K C�L��7�ſָ?���ݬ�a�T`���PX7��QE&s�o��,R��w*�7��y-t �}K*�x	��]�}�/�}��͂��Q{;;j�`�>H="�Vh�A�{*����b7aj{������}�!�g�ۃ�.+z�ת��I(*k��}�wl,,��e�rLq׎9H��DP m��j��\�@rh�Jɤn�H��X��������v'CE �A���P�X,�2`����d|�ėI����,��cG$Z�"ɏl�+w�����X텲���!�0�並��]�����,��W�V�ќ��>BZ�	2�=1.��؁�syp�ߝ\ �V����ɁT�����b�Ǒ��ZѩKλ�"��&^ʾr#�*����\܉`>J�+�`��
���%��v۸��u��Ӕ� �`On�K�s���a�J�iѤ�g�FF	 �u�!�])�ԃ����f�ap5����?�{�n�ʐ7�$"���՜�Ys�I\Q�w�+ݜG3y�	9���E��0� �o�:�.%e�� ��P+(Eu�RN����M5[Í����1�wo�7=�� �;�������D�Dz���b^2�����iڤ����S�%:��\��Y1g'�TCCo�~4����{|��V�W�:0�wB�{	�����ᖋ.�r� ��)�$ɨN�EX\�����d�}�쬬VU�N�@L���R:/����4`�j��ª=����}�,i��$���DEh��,UOM4t�J�n�=�qh�8��n�� '�����;ѩ����+`�+|��2ؤ�᯽H���}|"f���R��tu�<tg+-(غ�ز����������ԛP������+~����	��H��v��2�RuJ�<�5�9z��������MwH� Jz`�}��fm��1Z�=�����_X聑��+i�o*Z����v��q���z��6����2�\�c��l� aq���n䁄6�+����[$�ȋ`ؽ�l�U�]7K��vK�A6�so���(^�3��z���i�2�_��t1����O��-,� [� '��ݯoUl���Hi#���f���0������N�[�RN����o��G�cd$W.��c�-�A������6�lvRJ���(f�H�ƌo�<����V1A��7<c���x�S�j{c����W����
�D��}�v��i�\VN�m�wOh�2V��s��p�	�`����F���&���|a_�"�������vh pb���4_cS�f7�I	l*.�4�� ��YD0}�:��G!�W>��2R����s�+��G�n��.=j?�Ƽ;���Ƹ|�Ƙʷ�!i���C��M���A^��|��^?�K&*22�e�A�,��鄸�3j�;6�����|����ոƶ����
�i��	����l�m�k��3	�M����9���#3������y��h�@��M&�u����e��8يe���&��~M㔚].yR���--..>!2V%q?���\2X{�ˑЊm@^d|}}������:���! ��_)BȻ~�d�0&��ǜ�me����<�X�������/�c���{��&m����f�[��m9���_��#=��� ��p'k��������������|p�� ��2�#�X��]��#(�"&: |�u����Ɵ���WD����ܽ��` w�]��@x���q[�}�Q>y�����r�VRVZ����FL|�o��
+�.Xo�<�3Ü_��cz;�VLq��)���CI�oR~������1��qV��ԛ/>��.��d� t���	�K����������Y�Wc[��0�;���D�ڠ@yͣ���]e�3g��J,��st����������XX%�c��rU�K��U��������%p���mC���Ϯt�.-0;�B�#���Y^t��[Ob�� ��-���v�|n�N���O�H�]l��E	�y���[6�?_�7~��ӧi��ƅ��9f�}��њ���n��wH\V1�M#��FÐB�q��f~K�p��w����6嶳��W���@��OJ�������q���?o6wY�]r�q�T���f�'�t��8{\P�"��	�&;roX������ׯ_��,	$�H׺mw�2����oY��p�^+:�n��ѥ��0��"��9��|�r���A�Z3ʾ���?���h����mV���X1	7��/t
����䋙M�3ͮ�� wA^���o
>ظʝjjj���8�͛7'6�׿T���}��C���.�v���������}###�ִEY�o�}�,�7�,V!��ٙ�ޕ<y���ҝ�{��3|~�Y)o�[��(��ޓ�65o+,���3��ILy�i:r������#�������$�36�7���j�~A�c=�^�>��	\T��s[��h�NЖ�]akP{X-A�9�����֕��Ф�rԦIg�JǏ��j������^1iW�\5�n�?G�,I4�@Ru�ܐ����}����])�;f�o>�q�p�+-��H�����{�6��� �B�u����g�_|�D=gw o�~��6�#8Q]���fE�a ȩUJ��ˠ��T��ܦ�:��]������K��7�.�K��T�Z��-���;Q n�޽�U�YJ���0f�@�+��N¨W�jC�8��e�	q�8��:I\.s�Y��M�T��Y ㌕F�F/� }fE��*������{�y�n��}�6���KF�f������p�u;�`��H�
�f¥�{]�	��g�
���ڸ�?�݉
O��KA;g���h�#g[녹����c�^���p��)v?�ū)��MF�5�N��>�p�ˤs3o����B_�R�+߶�7���D�n� j[ #�?�i�D.�?���^�#ļ�� ����鼭�^�LK�O�Gˌ�tO"W�^-�@�	���QV��~#R,З_�����7��jV�A6>{�F`�{4�!���l?��#��S��y �~؏(��$/Bkw����41͠����T�i5^tw�#��_ k	Z���O>@������Ym����JFڒX���=
�|��� T������pv�\��'��$ebh�?�-�dsѸJ@�<6UGi�=��)~[⿹�(�r^D�OM}H6�OLL^{vы:Q$�3�����@����Gfw����{9~�9��E������\V��==mE�ĭV������Cn;M��ң)
?y{��nK�>r1�$���5���^�Ȳ����,��
��lpK�����=�(-}�y�P\/��q�z	js��u���CX�ddD���R����P�$V��E�~~~hb�������҉'N�RK��N��1��&��X�)���񰄄����7���o��F(lL����6�S�.�g͠���h��Y]�r�t}?Bl�8�l`��'���3���zBC�� d��~����g{mp�mw�mbT��²��Sڽ>�`D���مm(���0o;�^h���\�	�m#���0	���+��� �B�>�fu�S�Ý_�"P��SN�~8�z�R�?m��N]��B�D�b�������1� �'��6���p'���^"Q��y�3���Oj)�x����Q�����?�ni�)	�JtBZ��=
����O��)��Ԥ~ay{%/�yJ91@n�v3�9u�k̷o���՟�d��9����]��$���׮s	��k��������0�{	��\��;�(��p9�����X��h�}��K������YoZ�&8�ٵ��'f�q�v^���A��VׄMk�N<�W'f��]��'�P�!�IBb����X���l�dQp�֗I`���CU���'�*@�2;�TN���P�􌹏>l�	��(՛�C�F�@�r<�6��0���l�Q^AA!H!����x���8�W��(�[R�� ,��[���:`�X��Kcr=��nrg���"~�K@S[�?l��=&�$��j�ƪ� '<{pT w0b_�R�HPa��m<�RJ*�77�"{1��O-y�ب4��<�e���=�����G��$Z�4��������|�3�N�e�Iy�J�< R����J�1S\������E�=�S癝j̮,�C=���>��X�)���ի�;��>c��q;@+׬����Z	J���)pf}���3��Pbן��V|V;��B��yC��pT4���$.t"�.@�Xr\}z������B�n������f���<�Gb��˥JKw���t�=����c1xóKof,��,���[���]i��	�$�'eM�C�^W\�~{H��y�ξ)\h�� M�>��p�8�h�ߡ�T/�ʕ��b6������#��ݤ:�O�2Ra��3
�ɼz��*���בW^����L��/���|귐Co`/<cDt KO:��A�j�o][DD$��<�q'`ty�J�tϞ=[�~l'U+#���Ɠ����� +k�`y* ��ܹ����t�q)&I%�KM����w���Ed���H�i�C����@���q�_M���1%����=\�A�Z�L]:���F҇�y�Ը��@Ü�|1�� ��X۟7 �Mb���eYYB�^?˓X�%dvo���s1�����t�D�R��ǰv�9pK�C��8o�ttttd�ͳ���E}��������r�Z|;m���qAN�C��ܹs�s�� �ɵ�0���e<��9���T�Q��J�ڏ:^�v��UKɤWf���k6�e�!|��0N����B[O��䦦�Lu!%&&���8rk˪��HiQ���	d%����Ņ���g�$�f#e��B� $kA��'���8��.�F�y�����r1�u��,�2�e����j7�/��������7%�]�A�J6
�u�	��Pna[�uj<~88��/����:2�T������u@�Z���դ*�=9� I/		y���$l��j�������夔}#���#�hż}�9[�����P�&��/<$ㄬ�[}�. ��C��< tg.�3{/�tf.X����&�O����L���5���9ԧVX���-[[��+zk��"�w��0`��D7�����*0���c������.'�[���V���)��#�������b1���,c{9P	8?0��"�t������]�����js��d�2���L���W��fy�!�Do:�p��_>��x������)��3�S�"�A"��K"�*#�f����OET�Ӂ �ݺou�x�\'6�ω0�E��ř
Y�S'�/q��N9>o�YaV	�E�Wb���qK������<��}���NR���1�E���ន�J)ugI��O?��{3z ��IƟ���9%�O���G�Y���g�����N�@�;EEE�u�]�ȟ�\�2�����4U����k����5����r����*�=%T����s��OG�((v����"�j6I�{G���Y^�O��iJ��ɹ�_�UUU�{���܃D�S��1J;�)�l�	�7^�o��=^iV��6�uy�aB-.6A>�u �oQ�1_�>ݥ��+f��ʗr�"}
7Rj?U6�
������>H�"�f��h�)�~G�a�ϠwͷL�mmm�X�0X���k �!�|\�����A�5��8�X����bSҰ�y�5=�d��l����4D���9ORSVVvZ���Z�KGC:tXٸ_�lW�TIZ�rY��_5�E�l'��&)�	�+�>�؜�A�I�L�;z`��=�F�Wu����GO�3Gl�@�l_����#>~��%��K^���&��G$���J�֏F���7Y�37#83�:�R�D�P�z�[��8�eokhD����ߛ�DUK�p�z]��S�U'�i�9�9�]r�(��M����|��ڨ
����q10��+�ͭ� �q����� �r+pV/�O:A���ݵp�K�55�͏�c���[��xy�1����J�y+l���ƃrbE?,,LTF����1�n��'�g�N�o���&��Q�aM�� ��)J~~>^��pȝd�j�o߆=w�%)���6������Fr��@A��� ���p� ��s����=�=��"�~�EH���ت�5���N6���x�V�M�4)gN�VK)k37S�CS_ey��w��������J�3�fU�������'x��Ĩ���(X��ff �c@G����j�vX��s���EK��ٔ���%��LU~��/oѧ�P�>}��<�����6%p�{���n�����^UVV�?T��h�����E<���Y�̗1y���υ��_R�[j�z��� ĤG�,��t�[5V�2ۚ�S��MG	b���B5��;�,�iS}^Xb9EP�h��r�����#��[��YY���
H��p�~��r{���y� �=PQ<�!�-��b���Gv$�C9�����:3�~~sx����k����qصA��M!�P���_�4v6N�$����� S���y����	R4~!�6���O�s� NxEP0�M#-Y�����@ �&Z�W R�,Ļ�����N���Ч��6;�4A6�Y?B�d=�m���9��WK�V�`��ac��f��{z�ܲ�WL�'��X�5���.m�$&>�L������]��{��U =����MOW�o�b�H:�[�t��2�(
B#��Q�\����o�tr�2<��.��b��klMp��K��:_3�j]��������sT��T�P�
�+�2�o�@�	�Q�S�kRT�@*�as?}*,�>.�ZR��qq|�oo���W��L=��S����
����9���Pd����Wnϒ���㌃����݄�ޮ��͙S�@��KEzjs�Q�7A����P��r����u���AC��ۤ-G�RM�nKE�{{{#[߮����]B�����d�7�U�ђBxu(�5d4�������ީ�WfK�\��\ Uᠣ\ҿ�Ԭ<}�YwI)z}�3z)��A�\�ִ�∧������ȫۀ8��9a���@�ԑ#G��]�-�HN3�+l�1��a��Yɢ���O
�%�S��'P����*����vܬR��>٣L��������Uu�Ơ�k UZ��ű��������*�Ŕ�o%�d$<���&l��\{�I䂉��� V�|4�)�����UD�h{�^6���Q�{c�BE��֚S�KR���c����0��&5�\�)���p��� 5�H�����	�e��d/��Δ�����K�������ׯ�����e<��Ǌ>I�$Q�!|�0n�V�9���R��P����J�v��ap����� {��0j���;	��R����e2�
p<�f�����b �T��7o2{Xb��E�x���ȯ�	�����'''C0�:����Ѽ�/yc�1XNX��7�	��å��]lk_l�k�M���?h.�Z�&��k�y.?�;�>7Whddd�L�]EJuo܅��/�rVQ`�U�J�q��患`Т"Q�.��y���*��¹"�X���R�W�ڵ7/�/+���
%)%�^�О��l �Z�|1�l�Nɋ�k��\:�&�D4D�|ᛀ�� EO!?֣\/!Y��`����ޛ�A+�|���Q2���{��� �͊b77JB4�u���q�[
�L���5,�Q����ѳB.� ���9X���\�l�~ &�]P "%�:ݭ�����f��jUw���B,Y��S�����p�~\&�q��S L|�J����D���?*?�,5O�}�#�r����	��&�O���]����\�u�wΗ�D� ��0�}�L`/�R���5��\���l>"
`�'��ڲ-����9mm톞* [_(ɞ�.s������w 9�K�$��ê�`��]]]-|�6�
~� �['�`���B�4>nO��ѷ]Q(0	�l��1�] ��ޭOO��Bt�Fw��rwS��4g�M�v�u8��!�������Q�Q=u�������Rb2�
��<��2g��}��;J~�)_��K��I&����>}ը�P�{� ���}��	=pwy�������<�}���BX�ϣ<�!c�luz0<�����M�\4��j�����m�2�рZ��icХ���,'? ��=���|�a�R��%� �� JW�#�F��2=%/�}Z��A[�R�	
.�=�D�� hi��
"��`b��/��<����am��\������o� ���-i��r�a��y/����"c{PF�kg��J�t�������1ƅ3T���+W������F�%�]|vW^(�*������:L�)FYZJ���l�
G�Ϩݭ���!�#G���~�a��N����ɾ^�`,�G5���c^Ĥ�*xI$N��eBrr��W��+Y�f'�����O�T�-�!C67��)m�
1+U��5�V�#'��p���<�ĝ��￼�	���g��@��|ذ�e�X�,�����=D%~aSΣ!F��{��c�&�D=�.ǻB.��Y�:D�n�]����mQUᙨW�X,VϞ�9��ja�+�=\��F���Z�=�^� � �����.�f�^���oW�"���(�H����!��z2�i���;����A�z:���e'�����0/��'^Mr�[O�0�D�m�?��oI	��u?��P�9�oʿ17/۩��ș��˓<ɯ�����`����m��d�j]���M��z[�v r��E�0s�sdr8,z���N�O�N())����ea��Ӵ)��o��e��<V'��M/�������n����)X���u�>��xwCpp�$�2�wG�j �ߗ��$9�㲆uj(�,o����b�~K��t�'������_���_�F�V�X��\9�4?���ٳoD".��F�'���s���"7��&�"ke�_�$��Rz/Cco�ס�Ӏ�D���4�A��5��>�F�����-Q��e��wʹ(�4��*�s����������)�Ɣ��Z��%�Q��E3��O�寎�B��{=��J���f��n�B�2<<�~Wf�$M��N��_�^B�B���h�@��e�M�=fw�~���N�pI�˸��j���V,�!a
< �0��Kt��ܨ�jh_�s�}3ݶ��ʈsF��
��������`�i��
I=��]9))�o����*z.��Ʃ@g^� Q;�N��|��s^q113������õ3���\���
�:6��\�ZcԴ9����\$ I���Q���7�Y�9�ŗ^D)�7�������u�aoR��Z�Hx��$#�;F7����JEQhg!��R2�(��&�P��3�E��;WD���Q�������ǽ.Sw�<���94p��i���:�>&������)ۍ�f���������sx�{�S9xyyU��\f�2������"��+^e(br�i�Ə�+6�Ν���{b�A���h��1��V=�Coܭ5��Md��Hcso�
�S5U�_6��}.W����^��RY�uya!�"&�������k��4U����	6'SN�t��J�PL��}�׈s���J ��a==�����r gE�)�����r�dX�G��RSS���B��Uzh��{����8�ܶЯ��gE�\r�誡6�v&��t��ww*� ��TTU���ޤ�ޚ���� )p��o1�G�n��N��!�`!.�7X�ʘ������.pnE�z�p� 8�;��pS�9�"2���OaW�t-��1����ё��ml�ր�X^!ሴ���'K'�c��֮�蘨���drב2����"7R�ﺰ�<���4<c���3q��R�� �8���3BR���
�Ό�C^~�8B���ϱ��b��t=m�@k!�E�T�w/��GD`���.~skk��l]]ݣ���T�����
Q�4T/�\�� ~,ArR���/��5��￺��2$$�⚪E��'��P�:�%(�5m.י}z�X��?ueŹ�8�嶌���L���\<����$�2���)�=f|�_�.4���W�L�����Ȕ� \����`/᝛!� � >�����Bǽ�CJ� /Lu�_�{®/
��Ԗ����AB�rBc:X�Z�E�Ğm^0� �\�k��2����?�{��=R4��rv�V�v�v����
�5~�Gz�9(�ɰaj� Y��g����Nsq��xc�����L.�޳E�/�k*kJGf܌�������GxVԁ>�cm=�U��b�\mٛ�Z
yo��If�����$G�-��A���?W�,Q޵�й���q�[�/�Ģ�@��$Dr�!ނ�88(����|�k�CN��9�4�RJI�bB(���/�4X��C/���ΐ���NJ�i��މ{CQE��vN4��Wr<�c^^���@z��"��x��o�Bd��(��n���k
`U} � `�Bi��xB�2ov�	K��0,�K�uV[aeل#�����2������A(�������
�� S�7�F*����Ci���R&1F�^C�v�O'aŪ>�f�%6z _�}�}\�y9�h��P树c�A>���/���3��d�4��I_?�P��I�������Ѫ�WD���o��E���?���0�p�}_��μA�ee���=1�cb�?e>��N��A���8e[[�kk8���&g�^���Ÿ�--���")�����9���K�Wb���D_���>�k�
��Y�*��6K��/BŨ���Ul��y���-����e�Ҡ ��Ĉ��N��]��q����8ѿh�\n���f{��2�Qb�T��8��p��aQm���x<�9��Q$�� %*!i!RR"H*�(�Ѝr0@@�	��Z%�kah��y׳����]�˞��z⾟�r�*7�u^炼!S�&�x��\ȅ��^�h���']�>y�����;pA��Aw�v��y�W��3!�7���#R����VH��X�S�(��A�̃r�h�:�z���9����1�s|#���j�� ����S���^���w�d���NRHF�v�,O���=0�d�pX��?��c!�;�+�r��.��DU�J�g��ׇ�nS��S�B�=�V���Bugs؊��sK}n�r�ܮ��YCeVn�9!+�0��c\	�!K��+]��EX�=�%��?�X�y�"�
?������ON}q�ta>��X�E�)ro�h��<O�}m8��#�X2�sѨ�D����CR��ize�u��Y:˨)�a$H���G�,7�����/���&���W듉Q�{���p�٨�����ԯ_�~IP��{1 �B������ʾ�n���2�Wl�<(���l@pp0#�PT����W�,�/-��S�BȪ�!��k�Ry�1����jR^D�e�����-0�;��Î�]`pp�E��x��+�-�a�H5�4_D�Z�J0kߵ����p_Ӄ2���݄��թV9cZ��>}z7��?H1B����2'�NR�7�aȀ�����|D����b-#�D#�4�-xYE����2F���ǔ2"{�K��e5��RSb"S�3v^�j>��K�an�u�NN�޲@�#��ļ�ݗnnn6��C�>*�c�t�X^j�y�m#:����~��-�>E=ՠ��+�0-�y699�JqߡĽ!�j#(L�&Ѱ���wz� }�of�.�D=L\��t�Vg�3��������{9cg����N�j̥h��%mW�� ���QW�N������_�Kr������O�� ��60�8V!�x"c ���C�4w�D���6EK`����e��C:�8��g����cjb"���_Z�.�g�]~�Cc�����2��I���ꏏw-~���C�<xz�.��e�����+���M��%�@�firݟ
G�]����=�O�b¯���{�2W�56�9����F�KC{1"<܀�*��8�3�m"6���}��vR|�i��P��).;>ל���Ȋ��`�1�ѷ$�6{�B��pvUB�8M3�$�N!�5Y��`�3ΰ�S��f"��I|Qas)I��ιcէ�E� #�|��$+����y����|hN����gGR���m�q����Z}w|Z��lt�)3����#^a��ƎX��B@������wv2 '{�A�����x#��)�T�aD��-���R�D	�����❥�[Lݑ�~���ƨ�fHܿMy�|���;�N��a����Fp&�u"�2�H����η����`r4�^ԜN��jS�t�o�JI���u/��7��������
w���1) �'�ImI����J��yM<My��D�E����1����1*���!V��� BOa�,�>g
ٷS�9����Ã�e
�6R~�y��4e�,��θ��`G����P�hPHj�ߞ�o�(N�uXKK+.9��ltT�\X`�X p����iH�A�5jJǠ�W�����0�_%.��G�?�v�h��+z˞q��!�jd��C�$?�V6ZW]=ȧ���$�h}�N��������zc�!��h�Mc� ���_���]w�,�;>/�4�3p���v��a�1����p"}E��3�� qas!�iy�+�Dʾ���N%_S@��S�������,H7ŋ��i`	K������%�=<��yf�d���w<��=�����B�Z_��W�s6 `���V͍��o���[y�?X?�D/C������\��Q{ysrr4�����[��>wo�l��y���>�����x�|��Vʧ� �	�Y$�%l��n���Y���wZ����Wr1d��C��W��n��7�JǪf��XI����RGk򑹙���o�4��ۏ���A9���G����ꯅ�>�/04�|��]a-)��˓FrI*)C>�a���b�����=Y��UϿ&�J����!Q� E�=|>$ p����E� m�P�_K�	S��ѴS�C
��o#����x֭�O����V���4"n��:��9�ȉ���o��$5�fВ8�K�l�?I��:��������cn����Cz:/:�-�,q��Ŧ߱�,�g�tT��9�w�q��BNR�?L`�i��p��?;��?�k����sQ>�m�̧�f�bDh4�@pl���1#K����UJ������0D �KRR�!?1����䣼�[��I��M�<G�K��_����H'���ǂ\$�q����c����h�a���[�K0
�������pv��I"���4�"_�tf�JO-�K��޽"���jU���q���\�ӍCO�<���Sp��}��(�T�^^�Q���B�L Q�u��VR���}�jS����
\�����:�|�8��O>e@�]RX�rTD��%�cY��/F�Ҍ��;;k��^i�=������Z�m�A�����x�۷[ʥ{o�Z�g�U����c���N�k��rw�p��F�2��9�Cu�w�!��|:�W �%}� ,,<�A����S��X������bϧ�4��D�Ɣ�m���IGSq���*1�mmt�hY�9�����]r�g�+����B4� 0�w�E�7�m�\r���L7^��I?��Ő������Y]��T{�a;;v�����?�� HQ���-��PEB�|�I����t�awD�%���l
j\�;o�{�:9�3j��O/�5�i��5����u�Ij!�J$#�D��pƎ����8FĿ�������nݟI�_�b�m���_�KS{�_	����$`����O�*�c��ijff�4�;Tn��hF��C4�>=96u��(%b}�}E��|��: i���1�����u����r.��cPQQ��Ԥ���w��S��@8�6B�J"=�+&���T�ܞ���5M�.��v���9�(�G8Ą���q>�_�\���i�̔��1o��4XgM�-�bsv�ܷ� q�a�$��e}{�Zk����_���hCP�{�\՝M�F&��C��ʐݳ���:�mX5�܅k��B�R���p�/�����+��B���7~%�3ѨB�#�}y��ܦ[�E���?��.���^D�˰L`2}����wr�P�F��=t��nk#0�����
�dY��S5�&_�+G��V1,Bd������r�F��OHէ�L���3W���g�������P��S^ޥhוn��v�ֆ��G��� [o���?Ch����%H9�׍�����;�`vV	d��p8N��5�Il���K��y����__�&Z9mdI�}}��1�Gc�C�A�ED��+��a�^���K���6����s��G!�cb�*�@!/�a��x���0Բ1����_塤��~�`�۷kMأ��Kz���Ɨ�a�K�ME����"��G
(((xbl��&��ݑ�N��Z�]����c�+/��^��s!驫�������{�����y�=��u{����C�x_����CO���xbn�����/�a�5���7�%��L&��؍}�F�7Vɋ����&=���ZGmա���@���C �f��z�T�������"��Pw6����8�N�voG���<�d�\���́�6)�t�e_�m5L�[Y��i��ݦ,yR~z�i�D҇��53ǎ�(��'O���3���yO���%]V-?+	g&'�nl��NlGu=�}?��Lp�\����'��겲}W4S��*illAig=<�-��ұ�j��Yz��0h�e.�4^���_b�Hj��$.p,��႐M~�+�]u��c8�`DD�b���a���W�冐l����pÔ�#���CNWWw����Y�o�}��y$^���hRa�����!��j�S�)��,Qx�\Pݟ�Ԛ�i�^f&�����hiA��lE��yyy�Y�_��_����|���|�1�0��atoU#S_�v�M�	@����q�\Y0r����{ZHi/�'NW�}f�;�4hr&$��p5�����/�o���zF�D;pggܡOr ĝ*��>6�ot���I��D�$'׷����#Y9�}��Z�+��I=ܓ��E��v$C75塹��q��h�0�:l,���i��3�H@R����K{�����x�����'M�EV��K?�C�r��\������S�>p>��6��kaiy~�742�W?��Iϋ�r_���H�	�^f��r>���fw�g�_o�y*BZ�K���"_c�$�`Q�e)f�Gs�����E����B�G���^� fWd�h��@�N��L\�ƽ��8�/��sq�� ��Wl�@T��QY��:�/Y91;tHZ�JH<��QE�lh�Rbz��s5�S�2"W�a(D����Њ=�����w��X~ǜ#��%�:�	�?�_�j��I{���͕�j�^)F��&+�-L��q�?<_�S�|N%V# �곐un�FJy��u�0�<fEtܫ@v�]��x�3 �7�<i_�����&�7v!�a�EN*':�S�׶?{�<^y�1��1����Z�@+4ŋ/��8}���w�RH���I�?�/~LL����_��?��S.�5��Q��I
B�g�3��j����"rT+����t3����XS ����^�͵LLL0�	��<�1))^����1J"6G�"�����!�|e�X�������$�����ozr�&��S��Xv����Νu}�7W�K4�G�X��iG��y�8	��:i�f�B~�)XCW����f��q���HN�_�v
�Z�U�&��M/�l���D��'d���9��W|�r ��]'Q^h��N`�Y6�[�VW���e�ߵrl3�W��w�X)�ʀ���fǠ���䤡(��׋cM�)��1�{$�Q�m,�<�ۙ�}0
&x�d�vF����/7�c�s���U,�M��^��<%c?~��nѥ���Eg�Nl�1^�X����m=�W���T�G�����W���cYD�7>��:R(5_u4!XЛ5����첳1�� ��r��n�.�G���ȳvAD��K��G�Ù����c��cMx�{�, ���F<�0�]����?JR[Kq���ϝ߿��4�N���ܩ�oS|����������I�H�d9�xJ?8z�7@�@d0��Ť�	�H�Y&^�q-55��z#,��_���5-e7]�~X�nr�O�s�F�B���Z]cCuX��կe�//�Ox{��`�}dX!/u�y�ɀcj�HL,LL|�eJ?}
�)��0���������A�Rp/��D�4�����0/�浄�B���ƾ�|n5m>���O��ܨXB^͐C=����v��(�����.hb0ֈOߏ�+㒑��s��!��o���7�$ȒeI�bb�Y�9���?�}��l}���s,� ��=���;|�Y�L��^�����V�}���A�S�	ff�������L����l���Yq(3�{#�����+�'��)8+���m$�R�h�O���
v���0�(HsPg�3Q�w�C]�9����DUuY���r����yv+H�˨���{��v��-�"y�6K!88�ͦ� ���_��"�k���oZ^^�X�mq������?���Ø�ƠQ|��~Ǳ(Mmm�u�U�'O8G��v�Vٔ:yI�?�z�	������#�jwB���e9�of���-O%t����G|��iLg���"�s<�lE+--�Y�W����Ǐ��g�̴��E����bI���̴O����������c{���U8�V��m��EҴ��������e'�@���o��HnZ�!����{BQIo�����mb��i�LS��v6W�ns�Ϯ̌���e���0%u4y*�3�];����>b��>ڸ��|��Y����:π�^&E�4~W���0����~��x���0i�s�y��t_?3%����?q����'n�4���ܽ��<��b�4���<��>p+w��[��L��ݙr�ʄr��aU� W��եYِSTz�d�a�mΗD
yܧ~��%���Y[���*c_�/�� {6>5�}���#��	cЮ�-��L��x���a� ��qD�ܞ�roۅ.Ӌߓ̮����`���sX��e]|]�|?�s��mMK����D��RI��W������-S�%W�)��͎,"&��s��ᑏ��ė/_z	�B��G}�%oح�FG�)Z���y0�s�U'�F?�#��E���@�Q���qJf&�#ۖ���������݂ �p��D��R8���b�"=�������\n���7Zcj��o��5�W���.Y��R�Q�0�na��@"b	���B�&H����3���iK����h%f�Ǆ���0��ol�$�g3Yr'�n�;�x��p}�LwwvY� �#F� ϙ���]ڊ�fJ33+����qX-vTmH��@ˇ�g��kBYf$�y�cx�{��.R���hؗ"���1��٬7.3�2�L�� �Yɭ�5����v��wa�px�����r,�V�An�y�`itey�+�e��|̜�F檒:��u2��]�-?�JW�_���e��f�H���^�����z.k�8��gf�313Ϙ�QW��w[�ߔ�T7v'r7���䔌ߍʯ����'�|GB/ ���V{�'�Nܩ7�p�o���Q������
��V�]��f��J��0o-��0r���ቋ�TR���=~,��&���I�
o///γ'�YY}���<�_�|�B���,�!�")�-��\D�%�O�<�YxdUp>�j�\s(̰V�x�Zݦ�@k?[f��	��0���"�yH�E����I]��|������to3C��(�*�4��קB:��%�KZ<���ޘ��)��;�k��5����
;[�xb�awB����@@�"����L̡�-�u%%=��HT��Q��&�;��6p�444��ޙ(���P-5i��{��33��=	��o�m�<;q;�QB\��t�9,4� f�Ҿ@d~�{�D�T�" ʙ��H���GK�"���e&�<Y�B��/0��������^��E���ֶ�b�{E��K` "�,��LL�JpR#��'��lM_�-h�<3N��B[��zi{�x�/�>�{�&J�<6˦�A���%���[�m����a�����FBF�޽{�@�Jy�Y�����r���J��g�?�tC=]|����W���5ɋ!��bV-��j�Uw�ʊ��؆������4�p�H��t?�7\/kk��q�R]]�a XRD�.n-�/|Y]�����)�fY�|�Z�[g�+|���Ð��395%<�|�]�aK(���00
`�O��]���֮�%냇A]�y�(��m2��J��D������!-~����`y�n���=��0�TK����E��ա�B_�޶�4v�z���������[��v�J���=�C|j_2��7v���0	'eFn���1���T���]�fH/��eŴ)���r�׭��D�Qj~�����������lB�|N�$j�������"g}�YӃH&�W��q} �诸w�YdL,Z��Ai��h��M��H�<B�'��L�;��g�A����N�z�l����y�7c�����bzb�[�Q�U�-�J/k��C��yTd�������:�zy�ݏZ}�<�]{�� ?n�V���B��K�p�����I�+\ǣ�|@E���N9Kf��T4�7�Û�$ I�D�Ԩ�MH�m��9��r�#
_wuu���b�?����l���qd��&5���%ӡ�4��"�	U^�=��a^ի�a���1�Fc7$vK�h�q#�����eI&�ׇ��T����4�Μ��2����%2�!PxQv�v�B
%HC�5�����{[p����կ_�B#"�sJ#�%4l��j,�@7eq���3���i�͵/�.���^�>�i��9�>�FSa1P�0���V��,#�lV���z}�,F?:�Wb(uvv���C��ܩ^��_,#�E�l�5X��S=�i�%v���׭Sc�c����p�L����ț��tX�6��:M�azdz����i"��֔~�АA�O�j����_��CL:��F��@���uW��OV�e{[�G�k����^C��KWHK����<aeeu|��8��}��ϒ�g���]�&5��	��!ʾ�2�8~�ɏ�C�F��%c|5�eQ��2�޷ݸA��ŔC�~U�!7/W.��ZjllTt��^~䛁���[)�V��Agf5T�:�D&�dϞ=���_�gۥ��^�D\�N���[�tu62���-,F�x�ۙ12Q�k(�89;�''?��i�h���.lU2�����Э��݄d^�$��a/^�4ts���IxہTT\�yr���\�Z!��zn7��{�P�ҋ�!����U��/Nooo�~r�d��9�)3����O ���	�W��W�Tl/gZs��$<&���323� 9��_�8�d��̏trt g�'.��>7�G��+kn}^�3W�b��(!{S���p���r���Ϸ�v"6�����*2Bmmm�Xg¦�\����}/���ߍ[�4^��@� �X����0�27I7���D"���ˇ̈/Pԧ[byn�0�ܹ��E��^����92��x�")�gb�E��$:r1���!��Qg�K3j�஬��k�)����x� /RYcba�8�A��K2�;���ig4���KV1��&�����L�c#�ϻ~��>>hm�����Sd���YĬ%��
ku��~�AsZN{C��!�L9��Q�H��'&�ff��(��65%���N���z6�=��À��r��L��pስ����������c��,fg~<�O'�pɚ����ko��b��8����_P`w]_�k���ʞh��'�GpC��2��M<�߼bm4�&�O����LC�����.mic[��	/J��V�.���tV�r� ��3RRz�:��,��t�m�{3��Pچ馏?�c|�mT���xI���B�B��lu��_&F�*��7��\��f����U�ҭ�^�ɶd�'�IU"����_X�Wލog�q�����!�y1/�5���uJr}<ފ҇ӳ����(���y�}�(��y�/j>��qP�G�xD:��cJ��.k���u���������RTQ!elb"�d���]V���)fDc�G�@���e�� "�k<53�[WW�n]����J�����u��t��o�$�D���������q&����5��Qy�pdeG��n-�<�0$\q�ƙ+;lL(�3����={�J���j��/4]��v�>����E� �J_�����M�����|��0�������k��]d��P|j��u�������Z_b�w���{�9Z�{G\��K��`bKKY� wg�rI�=���mEn�ؤIi�^�K	�:QDL�-F��'y�g��]���l|�c�&t)���bWt�G����W
�7��ݹF���M�o7�}�uￕ�y�^+�W�H�0��r�ט&������p��i��V���3�x�&���>�B���~�����1�}�f�]�iV۟H� �wDƏ�5@�G�3g���L��>G[Y�D_-f�� ��\B���yq	f��5í��5��	��������c{��)�t�oH=J°�~c�b{�����bX-h),.΂ṇ� /��A?Rs�&{�p��;�V3oqW��tu�n����y v5�����l?+���g1�c�!�b�r"���$��hp΋/Xz�NPq�}$�ҍ�j���
IY���W�Yp��^#A"��E�������vg������n��(��?L�&�yK�\mck}�����9ώ�����\[������wWG3SIŁ��;�{pʢ-�c��Y[_����$�y��E����;Nߜ@0��g�_gJ���"YUC",���-C�k�*��T/t��x�>'cG��"�(��R�~4����SK$R:��⼛&�	��*����d�.XǮ����PRR��0�oIt`��25�p�ԃ4��t2v������;��}dwi	�'hiQ�i�{�d����zL��g����┙F=L��tU}�5�j�"$�����,�zp�.��L��}U���a��8�M%�_�g���oP6�)&��#�mhcs鱑�^�ܩV�-O���wX�:�s��*�x�5�-"v�-���XEӕ�PƋ\��]�7��c���-������@~g�ɝ�B��X�=�E)ȉ�H��|t[��5]}����3w^��cw�����I �HRprjᆈ�[h.+.u[��^cV؇�5i�"��.v4�;١�l��	�&����������׾Ͼ��:ވ��5��3��.���M��:��m^�hens���v��K�b�������}Q����bs\F��'8��I,�u�⿙�+6�f���%�M�]��u�i����+%�&��!�(>i�b�l�M���g7+�
�́��Y��G[��d���F�(���a�W�=�K�������Zbo%� <F�m1b��˗k�)K�KKK7�H��������<� I�.CSB),��k,��n�TW߅���F?�BR a��W�Z�4ƍ��IOZ�yk�q 漘�p^@f��;�*¢�8b.��&&&�� ��V�:�5��=���$��Y�k��mY�{�}Yw�
d%�O�z������H�"2�6�O�T���?��� �pޞܰEB���=+Fю�;���3�����*)����f�HI�W�����z�6�鸔'T��������C�F��Yq�c}�߱��Xc���S�\GW�-��H��� ��u��z��k#skd����ȩ�L'�RUuC���`n�@��'x�T+^��k��幩�Z�B����w�����|f8�^��ݟmmtC:�9ƫ�߄��S���e0u��1��.q��{`g�@21��L���	�̵âl����`,�?�~pt���.;/D�RR��O���x���ͽVU~���u���}�[��|bb���S��Z[OKԹ_�:�%�Xu����3(���2�;�L{xo����	yDX<~��f]|J�'��OW{�K���D�b��o���9Ӻ��U��@)��h�'��
���_���R��"���-˰��4�(��p
��h�8��ʯEGGG%����H!^Ӿ���%Z���?�^���̈́,]|f��s������h��u@��jp} �I次��	�tn��$G�꽑�����'��Į���B}��N��N�z)��Y���0=��eUm2���2R�lw5����iū���M8�)̍a�x�3ܚ]Z�T�qW]
?����Nd��9�O$-^�-Y���R�Z�a����#��]P@��	���{� ��u@�<����M�$���vX�ފ��i�Ȣ�ښ;_�>�_�d��-/67�§�E�}-|n�c��5P-�M��6����"���52UMf0�dꊕ�ϓ�IF���V���-t[3��#0��2�f�}eM��S'2���ҕ'���}�|��
�_E=�>�[hb�	f_��	Ȉ[Mwek��6�T�)J�+�k�����hG�~P}����I\a��=��2&��h�n��(5�V����j�e�a�������2w3q�*������X��_맔���ݷ��3N���z�׃���BB���φB���Xɥ�Α,g6dZ�g�oy���}�j�&DmU�y��c_e;���O�*8��e�����RfDs^L^&'��y�&)��ZT�rss�x��<�������<�+O��i���������{���ճ��q�����t*y��iqV�l3��;������}��91�U1տ$���������tzⁱ�T�	+�v6h����a��b�wQy�8�4u1���QF�o}뢨DHm]Ӿ���Z����|.�p�=���5i2��j~�LuXb�M�i���(�LNN�ef�7Q�o���������[T�A��l��� 8Ԫ$�{J�/��Q's7��L�T��4�N��
�y��lT�osoϦ�x2�"��ى�ncx�ZN��Pa�n�K�������P��K�՗�z ������]�}v��=��0�]�y�T���d6Up���P&|e���z�8�S��IB���O��8�>�-F��5O&IW�����a��38�3�����Q���'��@'v�`d+N�S��>��z�Kٻo�0d�!]�|��e:����?($*?���8��뗋����;J��6�"r*�ˈ���f=1�x�4jVۣ&�!��x۩,#�"�c��`8�j%���nooC��OvY��RŻ�n������ﯺ�4����x>}C�מ��wI��-�wp��9W���1J_N�TCRř��_b��*��Zv-���l)�C<үR/�-�~����\��x"��UMw''�BB�}��?�(��M+Euu�K�7�Ԯ/��;˷u:l�rR�����Q�������ܻ,/&J����]�t;�B�}��;��~iA����y���8�e����YP��2@j�099b7�L=UC3E!���gg����v�����
I�C��(�V֋�{��i��ӣf⬦�z��6M���)oN���Д�9*\�`N��a�N����?GiO#�- ,t|��oG/1܎���O�g�V���tAA�v)O�L�	�.���1�K�����-���\���c液֞�U��6/���j��Z�0�/]lü8+Ƽ�F����)տl��'�/��k���j8����{6y�,��g���a��@`_���ǆG���y<G�����t=3���]�a>hB.�-'����������1*Di#I

�R|6���`��B�I�~m橸��_�)t.�'iL�[��74�v���?��]MTv�I����y4F�!�
v�)p��biܶ�Y�u���6~44HsA���Ϗ���"R����6N|�܊�ASLS��eْ��K�#�����q:��#A����*�U�J��Ie���[�v�����hT��c7����\{`�W\����{�B=7FW[c��RSSU�N L( )�Kܕ�a�}O���fI�"��qC�ЕM�W���Ș~����S]�,ɒ"� ��0ו���0B�~�8-�+כ��^fA�Ί����C�Lq.�ݚ��X��p�TOeVDk���=��h#+�oPP��	�#r�z;OD4tՏ��l�P���J�u�#"�-���Ph⯩�v17�	-q�ԑʠ���=��Vo�	�mcf��=���M^,�]�.��
C�]��X�K���y���2�X"I��<�ѐ�Ԩy�[|[��#�K7�]�uh˅��?���{�ru�n�+4T���h����g���/#^7�m���|ԟ�.s���o���ގ=fb�xtR����uu1�(-e�	#��;�i$��������̞����:��x�幹$*�OX�(���N�iܝ����)�z�-g�*��I�T�@���?����\0���͜g~�K����L����cVV�&���;2֮3�|���
�ٟ����_�1��F�?�2r
���YBB�r�[��:�:����'��`0.fgs�8^z}2��D����֮�j�gB��	��3ŷZ�/�����S[-�O�a�ZؚX�:��wd48��&-	��RrV���(�܌*cYj*���v�`������܄Je�YP~i!��[�e�:��/�Px��
��;��k��G)���O�Q�7�*.�_^꿣`!�ƾg�K=����(�^"T��z$��+i�aqk;z�N������:��χ�C�N_�;���pU�ďzzz��l=62����wm-��:�K��L��`���Qt�S�ЬA��ן1_f���g���Xn�pK��kS\i�Y�V4�M��)I�%8�ʚ���z�)�A�2����ll����e}P��[@&֏M�	p�9XmD��f@��I<l�`�T�iIߵ<.�$�*��oπ	�pyr9�dj*^Dr�/�+�z��'�3�y�iS�bׇBj��Bu���ɻG�RD4�_����ܯ�/��lBϩ��E���.B�m�ۻSV+��wAy�3���U�ˢzr[W��(��)iohy�)�����O[9�%�f����6�_���WU��V��V���`�����/S�^������;~8�sO�Y�)Y�L��c���}l��<|�d/�4�c�aF�S���� Ȫr���Om�<���:؛N�ZD�T?1ڶ�5`�z��p9k���G[uuɏ�&)����A��O����3'e��s�N���r��b�rݸ\jO+��<���yaX��U��5�N�j1�?��{�����Pė���c �6%���Q�w�O��8ߡmQo$�0,;;��n�`M���Jy㘆��WJ�W���W��ʊs.���跏T��������/��g��K�\`M��J8�62,g�����gO��Ċ1]Ǭ���@A%�ڠ/#�	�|IM�c�����EW��r�y��`5��E�+�������c�XS��y8�X<f{)ISW�WU���r�x�C	�q�.��8�U�q7ļ�S~ךEJF�+o�LᎻ��,w���з՗��d����?�vݿ��q�Nnv|���eummf��k^��F�V�Y���� �XS���pb�Y/}@@�c��I܈��Z��1�]��S3r�}}���nOE��"�
�W�!�gyc��4>s_�\��ޓ|��Q����δ����Von���DAVSS��ѱ��J=Փ��֠X�(Qup��jKV�������IWWW��C<��OC�Dj����������ƔM������36y�.��{��B���"��7˰W��h>�۾��}(5�w��~���mm熦�?(��]چ+
��:Y�]ϞC��ty)E�J@\�%�_ׁd�lDbo޼i��)�M�#$~V�a��`�,"%M�I��i��1��NJL<��Sc�J_��5��rW�e�f�
JJ�]]�uy?��M�n�)..���Z^Z�㑜�����J(����G���F�<g�{��������Aq��~6��2��[�R�3��UG�n��C����˱㰂x��q�����s���	o]c%�W\Ӱ���/���߽{9vh5�����]��z���~�G�aw��7W4����ٞ�ak������KV�xu�r��K6G�a
f�꺚�8��A��Ll�$l���Wde}=�&����H���u���ך񑋋8�ѭ���K����]qN��\�\��� �/��zX�BX�ͻS2�����������2(e��8�gm��������un���E\V-^�j�\r�X�8�ڞ{)�S����"$B���R�}���	��-_����XnS��	meo�d�X�EُZ-��V��w�!MC\)b�Dz�ۃ��cE�׹T��ve�g�I'�j8QO�^w��>�fe�]�j��8��m�k@S�8�����hd؉]�L]�Ҋ��P��Evʴ�_&��		��G[�Y�^E����������
z}bQ�x>�&�.�>}���=��9��bu�V�Q*���d�枒�#:d����A�-4:�o~~>��(����3���� �	�t���&��`N�x���KmB
u�}gP�A������mm��אkB��F\I��	C���5`�냨��Q��oMn+����M������i))眜�a�Z	����,R��yy:��-:�ugc~���sF�y�.<�ؗ�Yk�8B�I���>oBLm�{�.<�!y�_�222宂-��gff.wEG�7e�S�I�ì�/�v�5ix�9>��4���������ś�oogw�v�]?\��
�K�A��J=��R���U���5D��[��J���������� ~J'�VR\WP���Ӹ��{���x*�ŭ� ��p�*Ű���t������Оkkk1�⡝���'����.��W���� K���>�� ���6&'��R��\���U6�46 U^$��C9.H^��3���wL(q�/��F3���_��*N
����>�<f��~��������رcˑ����L?�E��zg�b:'��i[�cwߴ���]�캱J�G;�w%�"����R�R���VqJ���TZ��	�
�[	}�������I�z�J$��þ<^�we�c���+t�LV ��0(��^��5~~����g4wt{� �pzȲ��3#?����WBܼ`� [O�N�"��g��R+]�Oq]�I�ȸ)�<�7�Lf�S2#S�D���@����U�����(U�t:���OT`�(�����le�s2q�/(�����vl���6����1`x���m�uu�<����O�m�l'�4��S�@ ���������$T�7�"	���_Na@$�i�V�����R?��
R$B���v�+���<���)��>���,6������Ϟ�V?�.=��(��'O������\\� U����K!��v��ѳޢ��1D��e�JPL1�)!X�d���g/B.C!c�Ö��NX� ��A�l�Z��R�ĕ�K���נ�5'��W[���-J�c
�X`��;7�AB��Ԟ>���@���JS�f@�e�(}Xi�٦<��Ȇ�*s����|B!TaTD4�2\�?V�d��ֶ��SB�x�n�򤪦D~V�}gu��WS���a蟀�'�`W�-(v#)ƍ�}s�����H�|IXx,kci�f��������jj�ƦJ3؟����.̂��:@����/(
4��9��$S�.�1�F�ޞ����~_dk2tK�]_��'vP1'̎��b?"Q��8�1��j?s�x��Ζ.=5��P
��%v�E��+�V044�1�`��c�A��5~�����>???�	�W�ۙ�mʗɉҍ��&l��	��('�� �b����k�Ւ�Hu��LU#���%�=�n^�t�-LL��<�y�ᱼ�<(�V���!�n��|���%��b�j\�p$#�����rs/B�y�������"���y�ig�	( (�)���ȴ1"Y~���%g�L���Dx����R	-�Zg�z$r����M;kR����'G�}�,�|�<<<�X(3��E��3��+KE
��s��_}�|��H�s	@b��I�ݹF����޲В@�,�����T\슦ׄ�l��a\�%*�|Fw��`L5TG�C�@(�/o5�<?��w	A~��Snb�{'�c`~��q�Q��QBN΅B��V�C�"n��DO4a�������nL�"�F��]��� GԆ�@�-�Ȝ�n( ��������!?��JC��a�a��K����Ǐ9
���C���&--}IPP�=�5��1X-ūxl׊��I�L��n��J#��x{�QQ���"�B��誏�!Ľp�'\�G������R���)�O���Ϯ�Qs�IU�'宎:�~�Rl0��corv.b#�m�1��>>��]q���~V������-�!K:�U;�P�
��312�b�w�W��*Fo��[N�d[I_:˘��s)5�H�$��O��}�n�Pb�\2��;3@�/+N�]�\7�IJ5��W�� �)��������"�<.)!�{�w����O,,��bѥP�7�����A�7��8l��1��c����2`:J�XP��ed	����X`^��~�0����Z�ET�������HI��(�|kS�����^uuuB��=	��.4%HW�>U��,S/m�0�&�B� �-�\�i$���UWW#���:1l��$�"$ߎ���9�aA�����+����l��!�3OGB�t�TT��M����[�IIg1��^���s��?~� ��������k|Ho���Y[k�O����%�{G�w��sqY)�Ç_&�t~��מ&�??�����vr��2�I֛t~���o&&&�w8�hv!�����V�R��S�Es-�+���,NKO�4��}�0;��K�A�---�[�j��'B��F��Ȃ�Gl�b^C���K�+�G6��"�~�"�vOtGn6�#Ey��Wv�/�'8'����M�ܜ%����
�����#�>�`ga��M�`c��X�x��/&d4�{&��n�^k��1}.��M��yަ)Hz�XV.��]��JV��J���3�UU�0,
�)n�I?lP���������yŧb�H@��FR�x�.��
hT��o���x�k:z�
�ܒ����+F�}k�;���=��3k�e�(M�럩?�?���M����y���4�#̪'Z�r��/|�w�hn��K�����������?v��vݼq��"��?Ӛ�x-���[���������l������b�d��ƿ?�ܽ;Y�lwO�I���b_��}�3��T��T/����#]��9E�[Ь'P��eW�l�߼��9s�A�~��Ck�8��|��_Й�ӗ.���G�jֻ�F�^O-��?��,��{��HxQP�� �,@%�DP�[JjAbW�,�@Q��\`iD��ea���������}f�s�{�w��̚7�����M�)�Rr=����6.<7/�:��ꚇa��<U���R#|��D7c�(;���O+�~E^xyE�_9���m�k89X>O�{�M��[�Q��<<����ן;s��+d_���b��*
����~�m]�F-�C5kݧ��CB6�9Iڬ�~��&�.zr�A��z��R��:�^�?��L��ϝ��0���=a�*�e7�fs�[�C�	�������<y��β����g���~������v��1�⧼�EW�us[��0E�U+���1Զ]��]��܆��q@<�b�3�9+�ЕK�s	+{�u���Km35144]	��[��:辌���;H��v�RО:�>�L.������uq'���X�����{,-,
���;�\	A�ijژ[�1���#���?��\��W�E=ߦp�6���57@�*��Q�)�J�r���UE��>�׻gV��Rbb*J��4ȥB��wJ��?�	���X���Cz�~ӡ-�e���PX�t�v��w���2�M�]3#�;���v�T�����X��2�M���j.jgA`�t)��e�B
.&5��t��y��@��T�^6K~[;Ron�q�{�٧�HV=K��w�����/�ʵ5�����z{�.B���Nj��#�� �Z_@z+#V�Y�͉LS�Fr"�w3p��u�)��˵*���A���L�$#��Ø�(�f���w\����ѫ3;t�at��G��)������1�Ce�x�:��ê��6e�h�*+n������u����#�(4L�F��*��dO��`H�˭�4'���{mo~O-�1�$%�Oѩ��/_����p����G��L��#i���-���~����6���ז#�$��l�[y�+�b��ݟ�3������s��߈0���G
b�D�����I^Ф�����p.\��4�Q��R�H�0��sr
i)u�F� ����q�Į�(�h���{���@lM� :#��V�QH3v��9i@µB~7����7?٬N���+O�(5�wZ�e��/bD:����ب��OZA{]�9�2���i�}j�i��:��@Ћ�nf��WW���p�{�M%��Ӂ&�2� A�fgg�n�ƽ�W"[XZQ��iX���H�'P��`S�3%%��֭�%���.=�{�u�V^��� �I:��'4��J��}m�n�w07n���!���Owf����D������:m��n]���&��9�q<�LJJ���{��K���t{��)p�ZL ��wb�'���]�.�#]h��'�޽{!��x�k���B3�ϒ�%�i}T���1,=��{1����[0����h,��So�9#9R��.��@�hӜ�S_���2�%&f7�)��@)�_�h�n�S����[46�={�N���wFV7�k�G�N5�)(�ЙZz���P[z8G
��wm�勿���JA�s
Mo�/紻AjR�(2Xo
�}%��Ҷ���Mռ�lMJ��9�M/�wR�"ݧG�˼R�7^A%'<w��ںʍx�*fɎ����J^��!+�*�Y���H�R��z�K��ZrcO7oΊ� Q�b�#��%��I��Zg%[����^�&Օr��ĊJ�96��C#M?���v�S��=ʷ_��gΞ���u�Ƹi||<�c��v��x_5���U[�ӱ��7Q���$P�i��)gb��Zn������~���ب�~�i_�$�y��G��݆�s�]��U��|�u�y��Dy��Q���#��"�!�]F8	�p�Xg�iU�#��Y��ϯN�Zz:?3�Y/S�����͛q�8��OeK(��M�l���$Gp.u͉��4O�8�Q9Eyɮ'!@9�)}�Bd�ޣ�fu�V�h�/m��bS��������_�Kݧ�'2S����{81��**��� ��o3q��2%p*���U$�"$d|)6�k�C���!��@py}߾}8���Cġ�h-����(�-� c�� ���#�yL����9����;�O��g	Y������[�U(,�,�I�_��	�&nq+Ǥ�5^��l�q����G��n�QW��J����H�gN��%�:W�܎�ZZ��������,�1}�aJ�����|
��Q�����
�������z�Q6ݍ7ZWӣ�f��括�LXI�X��	���d��<�)[~g�qN��?~?��H���J�"�_@<�7Ͷc)5��9���?�˗��f����L��8ȡϟ灞ck�� �ƽ��)�ѻy"�T�aR��Fu�3�SCM��^�},�OS�rѹ�3�����c@n*X�)j�w?�G��Ivþ�W�ߔ.��a����V6�2(X��Wqq�i��`7�+W�����SF>%qڱ�:H�ųb"���7>h˶���LN��;�;P
6���}�Cs���8�H�2"�a�9���׺��gǪ�r0Z�+�E׮7E+�����Q_�%B�TG�㠴4I�;��N���j:��*z�P�e=�d��\�䤕�v�������dM�i��1G���I:;r�ǂ�A3��:Ɂf<���Eyq�x{����%�Xە奰�.	Va�x�*���y1ۇ@a}@���+<�S�1����.v�~�;%�Љ�UtXS0g��%�J%����Ë���<yҝ���6�3#lɄ�'�u|����9�k:��_�9wn�:����8׷~������xAu�����Dp	))5�8���%2�,$�0ՏO�8�W�"�����`��OG�'���DW1��f��}��Q����g>�rv��䒃P:Zo�7K�j�e���;�jjkW����5���x%�ׁGD'k^�"��c���6�b�}�cM���� �-eGɍ����,�8��~�37�u�2P�+:Fn�ђ+�9��ǜ�E|���FB����F^ޯ�lm�:!���G��A�!(���Y�M�{wf��h��謰� z<W�ŁZܚ��*�2J�T�:ݯ! ��~�.x}U� #�1��@����E��+Q,io~t��}>�r1�x�%�l�8x�(K��U�@1(�,�����>L�h���%L���ưx~j��ףU��:��ܵ�<e�%�����G:�a����	>+��ā�J����ð^ 4�"\̢�6�];���x�葓�nB�.���!�����%���7�=���#�1�M��蝠C��9}�d���5��e��`χ����U�
{� o)2�dh�x�fQ������&t?:�i6.�󘱙Yl�ϊ�ׯ�bn�'�C�[\IÅE?�JW��ɑ�l�����h^c=�Z��z{e������c��ʋ�.[�һC���K�f�ڟK� i�/�E�C��mȑ�i���<�B���|N��]v��v:'O�`ê6�o���%�o�����yA"������*+s��}��	���!Uq!? 3�������[G��I�����s&U��:o�D":�\iM�ni�¿�p$���0vUݜ˕��C��r����eF��N}�<f���q���C�}�XD̗���d������H'�V���[@��E��ۏ钭���F�
O��c$(9��>�FYT+'x٫�*�?[�N�q�tl?�zs�G�Ǐ�>��!b�����tW�i���kx����Xi�*$ucFՎ>����.�r��gˈ\��ֶs��oQr��]��N���բP�,pf3%%�� �.V��~�I� ��3`<k%7���d8rH���<
:3)1
Då�c+88{����aȬ�̳kP�$�]+D<�R�F�:�,�AF�0.!�$�G�ɚ�n��]$G���ȕ����#�.F+�*�˦͂Sr�� ��?z�1�,=,���,&����榨��o\� k����V�d�����5�
��ND�Q�'J�Kb���2&VuKVwy*�G����RHɠ(W���n��m�v�IYd#^Ne|��Q�SL⠜�T˨�/��ʀ��p�t�v���l� ��܄V�"��F��2��;D0�t�O^o��-/7PYC�8���ù���U��j��Tַ?l;�̊����z��V]&�Pi���f��E 7v��|\yfR���R����ZZ]���(s���_BW^V���W{Jn���[��� �]>Ho�� _db�reم�|϶�_`�RA��׷�l�mW�,{�����>����vD��v�:��F0�[n\M���燿���c�7=v�o!_�؃q�C/п/66���z�gϞ�B/�T�lU��W�ib�c�QH���	)��7��3C��1�=hP[�����ر���u[�f����)�9�����4'�6�����7O�R��iG�3�W�e���K�� &y2�aĮ&-�k$3�;[4��Z
Vw��<����6����c\�m��,�����9�P��Ƭ 8Ȉp0�bd�L��1�i[��ٯ�v�J� !��s�^�0HM��/w��^�@	����J��o��I1;���7�@�l���2iN�y�p��'����zi���È��4�R��[>ǝfqj��R��}�5�(��)�-�sH���1�bW��-��=��)]ɉ�Ym�������T��Р�(��4�v���%C���ɔ,kwLu��ݻ��9~~察o�c����0[Qyy�V>E)y0�(v��՟�ݿ�kRF��;IzV i�h���TT�Yg Su		;���.�d��EQ$���*{J=�����rJ܂G�1��i�{{��m6��7������eu`ڵkW2� \�Ms��j%�ZY����KXU���W<_���S�B��^��M��.PF����ə�#n�LD��W>K�>6���C�Ee(X
�.=�jJ22�sssGn�ǀ[{)��~��;n#4f�mn� 2V0ߖ;:"7�M�1�=�+�~�<ƬL.��o7nN�Z+H(<|cfB`t <}Ɣ��|��QsQ4XP��!
aN�!�6Ns�	���	ݼlH+��iJ���r��A�L�&~�x]Ĉ���e�/�rb��(7��v4��|��5j�G�޾}�Ht��G�,ZO�Rt���;dD4�;������^���sf � �תu��_:�2��̈v�T��h�;vTsrSR��=z��#/����9�st���K��XM�{�q�/o��o�X҄0'�i�#����۶��ϵ��N���� : R�oNX1T����CT�}��>�r�PV������`b�~�{���?�I��}ۏ�S螧����ϻ��z��\�M ��?R�MV}.&9"�bl$M�l�J�n����--���#\�.�K�H�Y���`
��}����D�s�b��rr�����Ͼ���d�dC�<?ƌ���BD/F$�۵���z˼��M�_g��w;ݢ<Z��c�&5����箂���9����55vvv܋_e�9�jR�X6��H*nb YN�����������]����w��-5�,��Jp,�j����rXd�]������Q%R�K?׺��&H`*7z������z�y�m!�}��0"# ��;*R�V󑳄�Xq�.'9������JK0e�N�~��dՔ�)&/�t
�Xۦ���њ�3~�H<oI:*	 �]4�AIB`�0(����Aݰ����|D���D����m�k8��\� ��	�"�wI_�q�cz����]g�G�	�`�S�o��œh��R!�
��m�+�b���;-�zJ�_�|A+�׾#�2��R̎�0 H��A�M���A��`�b`���F'�ͪ��?��|�1J��i	5�N&Ӌ�H��8�u�r���6q������p)1�}X�˜8u��3<%\�M�q�Y}�j|8�[��	��|n�\`��b7G�gl����k֡l���,���9�����Y1�m4����J�_��+Sn��������ɨ|w�S�-4C����hQ*(�|��N�S��s=6ꖎ��R���?B�� |c"��8s�-,��d�QĊ���hۺ���߸0����������&��U i�*݇�Iy�K��{{�fEy�:���y̓��;�[��_�.��s[`�@΢!t^��P�Z�>��CW^1ͲG�!'LM@�06�}��C<����>\ H��-V1f~и��miz;�q~�\�<եQ	p�?�eW�>�Y��rsi�����y���a����kMH%����"l��q�ʕ��U�C s��z�L��I��e�8H�Ȗ���RRe�0ܖYX6gŁ�6� 6�
�Ϳ����+��W4))�Fs|������Y��T�j������.՛��]**&�*˅��%��X�j����gaaQ�g�0ć�-� y�S�/���/���rp��v�`��@2��$$%�6R��z�G����24G���̎��Ǉ��EA.U՟�q]ygѭ��f:���^����Ϯ����H���� ���^ЦҤlt�SdV�k6��+�S���~���y:X�MǗ�P�F�m.����K����%x��nۙ�("i�J�3K�=�(�q"�0{�*}Jz� ��Z�0���tQ���=\�L�!�JБ'���t����n�k�S�fz������^cg��X�ii|�LU�1}{Lcg^��$���Q*6��桎���f���c����f1ɧ����Q�efu�"b�Q#�H���G�O6O��7�6ґM�Q�fѕ_���m��P�X�$�v饱��L2>U3qU�t�8�A��^�s�%29ʄ�=g�ǩ:w�����T[�@��u����}�6�˗[Jn� kC��BO<`�w��dQ�]��t�V,��,��+�k�`��\1m�L��g�f�x.�gvZG��Œ�2��H��{C=�A�A��5�KN�ƢjP1�mG��-9��r(��7��L�+~Jp�S����rO~6���䤫��U�~�؄�V��\��í�1�T��A~�O�Ln�Q�,&��>�3��.��Mc�#�ɢ2IB�����~���,���V9T6]���;����ׯ������mZ��7E[��!*�󓹧���e�����Ǐq.ma�u�]-���K�G箄6|�n����wT=�5fY*�f���^�\f�E`�j�p�I����oI����,ы����2ߓ|Ӵ ��53�h��j���bt���89Ѳ�fN�>wl,��J�X����mmU�X7�l�}gSÄ��9�*Q2�XڨUTT�H�0ߕ��=F�!��$$��΀���������۔ǖ��$� hUt�A����H�&jRC�/'_#=h"�k�	bԚi|�#�3�R�xy�Hx��BG[;��4z�`i�$�� 7�n3����Y�����ܤF�m}���<m�3��羇RK��cϨW��4����v��ZВv�����.��[6��Jk)-�����lG�-=i�{�i�rq>�]��=%z�	����_M�Id�>�Y��c+�E������I�^b9�:m�ضu���Ʀӌ��Y:JS�����O�-�x���)֕�� ǭȸ8p�*!�^�A�R�ӥ�mhI��M�����J���g��a�s���V�rN��ܥp%�Ps���Z	�թ5je���Osت���b%b̎���T�bYJ!ς�^3y��g�P�?���y[X���&E�um�t��sg�^rw/&V�u�g��n��H ��2&����$醗�t���� 8�"6���v9�O�[d�#��z����]y6_�[ߊF;Hv�ĩ}d�t��G;/�?�r��0�mC��80�K�Q�f�N����q��cO0�\�h������
ge����O��Y�v+$3���Ef�����5j@��^���s���![�rl���� ��H�Z�ꙗ�痻bHt��iFb���G�B����V�aR�pq�ܭO��Moe���$$$�dei`ef���[�|Y�4R��W�U+��}��]������H��$�I�`O�y�C�~�����L���{d��p.F����~hvS]�j��(и�xt*�s8J�ѡ�.�m���"�v�E�K���A���ٟ_�._��_ 4�#ܱx��QR�G��Dۯd������=��P%�)��'�@��>�aM���m����@����i������#��j�Z��ٸ�6M�kV8�B�=+2-)�/��8�H��AuyQ�͙��ie���Gp)�)�o�!�ɇ]Ա��0�9��1Qژ��6����3����2��84]�D��]&�F[d�4V��8]�K4 c���6�f���y�㤍,�5���_�2)3��^r+��hW��f���(�������hG������vL`�DnMU��1:5�?n]A��
+s��4��ALE�/�3���:��ބ�-�tF+�qf�.�")r�="d"p�~M��u����Xڝ�S�Y,[i���"�PN�zs��ut@�;#>o���i,�,~�R|��Y��G��欢�Ү��ӗK7=�����N����b4����Eϥ�F�6����bҷa�/�X���ێ}�l��{�U��z��bA}�釫U�3�_W7|V��U�T��]�
�M��@K�S��k�6�	ED�S��I�Q�~��'O~E2�������+�	���`�il�&���\�ZLNnnk��z�m���T�d%��[�X�BI�;&�?lB����E�y>+�ۜ����w9tPj��Ѓ²vmͦ'��{R�5'��2!�n�w��M��P$Î_/��̪��&''K����d�7����~�wx�1��F�NӍ�I%�z����ۻ*�T��cT�_/}��8�#;�~?��AA���}E��D��;/�A��0OV�ȇ�����Ţ]�]��ojIP�%���;d��u��+��̴/m�&���^�܊�ī���ȍ4��|n��V��ǦhO���ٞ#��{7'�Ǳ������M�����n �W��-P�j�<����ߔ�t�=3��-���b�`R�p��[yV�����4.�u,_�3�TɎ)��LO���V~����gX]��aG�J����r��B�M�Lk;ШX���V�Z�1����s��G!�I�8���Y]%]s{�����+\�'m�7�	{��ǰh��ȟ�< Δ�<�ӳ�Ϗqՙ˗(�E�%1U��8_:����-:{DΚu�h���NWg/wZ�Sm �?�������]bb�,jz����^SZYG� g^�-�B�D�ze����#?q�:PUR=�b�������kf5ܖ�<ׯel,=�Ba�ښ$���<�-e�|k�ǣ����/2w��X��M�Ne,�%���6$���gy�� 
�畎Wq��0�^�:���u�q�����P�6�c?��nJf�5�5mظq��g!��(11��w}���Z�cg7֚
>��ܻ+X�ΥK�:�7O���E׃���7������d�+�NwE�?^^�˗aŤ��%�F�V�|a��o�ز�A]i*d-Ko~�����I����^��es	����9Tg����_?k�%��j�h�3�}���o�=����,��۷W����S%�|k)�U�y�ͷi>��ǡ��2�>���X�&V�+@��~��\����$��C�A���Nl2;����~>�$<;��tO"C��5o���N$ c�6;^�M>)��7s0�t���w�+���m���
q�(���e[�($u,�q�#Z��6�=�>y��M��ۗ�1zp��D���K�s�-=\a��G�D<C�j��wy�&�]����d�D�uX�tNX=w#���n�ʞ�z6"�<��.m��3���0�DT�y���"�x-:��|��m���h�-��g:�:Q�����^�Q	MD`�ɏ���Ցef��!�QV�W�[W_�,�?g�*�yu��t�ɞ={n����+PM����'��0�f���[M�Ӥ��ϙ��S�Z���@��a�Sz�-�fzdľ*i%pɘִ!�ڛ:V�/�;�}��.j�W���� 3D%���=y�4G�Ӱ�!!����x��@�Hg����ލZ����^f�%Yӏ�s׮A �W����b���R�	
�,f׋.�~v�,��ޅ)<6=�j�!��P�4廝���r���Jb=Z�����s���e�uj՜�v�R�n-3h�L_&�o��6�9k��ts���!�:�t[<j'��:��Ai�Á=��b��]B�#j�yH��5[�S���>�^����z��'?׼��t��}�Qd��c�b����g�V�����e�?F����T�^OM��n���m>A�C���� [�y,��Al���$����QɄ����L�)��oް��Ȇ�(�K�R�S1���	��3.d��ZU��K�#*Д$t2��ۧ�u6)�}k�Ru����[oo1n|���d�h{���}��^��ɦ��4_�h;��Ok�c�2���ϯ��]����ɺ1�X���~���'�u���S�����?��
d�~���K�5�5'��#W�l�$ b�����^3�Z��{������8���v!I�>��?R���BX��UAkh_;�Ny��* �y��Ξ;ׄ����z���3$	�]���f�̿4����E =&.��O�E�ض�0u
�V ��.A�
��ˏ=��R�=����rO=�[Xx�R��z�]S�e��қ?v>�w<`ݿ"��ٽ����R��/Wc�z�
տ�u���V^�`�����G��x�̒˘� |0[�ކ�F!C�eDP��l�  �OH������C��F*sߞq�5\ U6{O���4�����l��?6�����S1rf.�?��8d.���s'\~|X�"�LP�:�ӿ،�RR�Ӗ��v��w�ܻt�O	ӟ�AP h	P�}˅pg������2ҙ{�>F?|�0}Aw�Ne9���][����p&Y�����>#<�r���j����q`���v���u�JMKk��y��!�����p\�{�vα�,�
R�����O�پ��#6e��f�wM<�Ժr���Z�H��}�+4��*�����s�`�����S/X���k[�7oN>zkͥ��{��ׇZv����|2'']ؤQ'���;�Z�
A��M|���KR���t���Q�`�<�������ّ�w���ĭ֙���ڶ�7oN0�	A���{�k7����[�>��i�@Jj���A�g�޻w�yś����mz}�x�N�GNo?�k��>����V�����OZY���H�('
��sQ��K��f��DF�<뫺z���� ��ċ~+�̇�L�u_l%c#��ԉ�7u��u���F~~���;N���<F=����6���Xl�"�vc@�+NJ����b���v]yɸ�)myUZo-s7�J�>�������z�M��Q�)�}�2�}�ϯ�qesV�_��I��������
k��!��dw*��]��즅�rC]`K�>lj�=��z�O\��c�9��4u'��~�N���D,�^�J+�A��E[�v�}t�j���9�5mx��3F�"CRa�.:"��G{;���}�ތ v0e���/f��%�����3�b�{$%7H�cJ/:��`0.S��6�����m��,ƈ�pE�����t�}3���v~]L�f��Ҳ�7���,͸���۪]�~>T�͑��H������X��V�!��e����̉ǘE��Kś9�&&�'Ο9�I���'���+��9l�2W��F���2���3-���y՘�]���=x�����lV���"c�G����s.l V M"R�\���F�����Z�����g#C""Ҫ�9TMo�P	�^�|/k��0���yN}���vSi��d-��l��)����lc�K����K�'l|U�uv��6'r�>~�F������1��^����`:��o�<�����؊�P���	+�����ܮ�ۿ�6X"��̋l��E,:M�1r�U�����g:ƗN��75R<�n���}�nʐ����-��J������n)��2�w����ɜ�����&��'�Y�J�5�	����~F�i�En����v�<���9�.��ށ@�"�/	���f�/�]����]k�3���!�p�=��)lY��/Y��+�?���x.0	�N�3�05�L��ߵI�T(h� j�o��Y���m$"L��\�(������s���Q��ӻDE�W`��T@�}<����� �> |��O��7&^i�������&y	�nw�*�@�<�~0V�B���_��ꞡ�T1l�$�)�0�+�i�w쨮|�xGk�i�m��v�,�k�U V����9�@�x��MAC��,�߳��D�W�]f�����ztBAdܾ�D�����nP�����)����>h��f�V��&� ��?���#�
�u���Gş�ϼ�Q.��ݻwKKh����|��]y�B���+| V��?��i����]~uI[�9��ț�t*�Eĩteya�#;D��ߞD]x���͛7�H���(8�`�;z�5��ue�>F������0[l�,�%���R��JY�ӥ�~�~��J�M�*v�EL��ǅ�ׯ3�톱&�)k��Du+�l��7"������=���i�Đ��<b�P�T�yy6�(Բo�K��*��z��}*CZ��7��/6+o�y�p�J�MUc�D�UX�؛1��c�
�� �Iǧ�k
V�+6�ަx�O�F�a�e�b�����L�pj�*�_f�th)ǝ��G:�ϝ=���˵"Y@��W`��)@�l^#�ti��遐R��Ǧ����S:�-`j��K�/@:��6�镶�u��q����0���f�Ȯ���C�qb� ���}D��Af�(�5D�����E55-3�X���e�����x%�����)�i� f���-'��W��l��v�r�|=Yo��d+�F ��C-�{����y�޴���*P��Q�W ��@a�$`9��M��f��x�@��g�U��)6\\j`�{��:zz/1�D7:s,Q�6ւDz0Z�I�N��OukG��؍�7�x<#�p]Y��aQ�^˺�T�$��Y��c����ͷ�yR��	X*f�ʮ_ް�E)��vҷ&�o[��U���7r/Q���m�\��3�U��~�s	��h��IZTt��;
y	����P-�8X�ȍ�=�[��5�W��O��n�����B�3��r�^Sv���k������7�m����1ô�л�P*^=9Qq��a�����K����L����d�1b=��
-Q:����2%ӏ�ד@�<����,~D�޷*6�vU�l�`Z�dD�	�#�a�՞��N"1Q�T�,����	̯Fz&z���u<��}>���,����dI�n��e����a�0�Nt�qv|�UC���Ƶ��iT���U�Jf�Xx(ݤ�`\��5����&{<��/[X���F�c���S���W��a~��݁�Ȣ�q�ˉ�PT���� V���U��M\ ��,rH����?�c�bi�A������� ��l6�|���
�ʪ㺐��}��U�72�h�q�si�-��t��DV[��с�qJո���Q�4**::���42b��S�& 0�p$����4e  ��ac��n<V+C���A�w*��1I����)��[JA�� �����ܣ�u�_�y-��<���|бGqi�ʟf���\^���ܴW�Z���$-j�:��\�TT�	]UH9�ݰ�D����ԣ�7��_�-$I��K~4FgF)y�X�?g�)��y���ޡ^�Er�L�(>W1�STt���)��X�Cc��|��J2���%%o�о�`-!݀ԆD��;l�w����I=���Ek�P?�nʏ�ta�k��c�&�'�o��>=f1�S��ӍΆ�æj�~���ֻ0V2����6���LuWT��L]��w�t��x�B,�:���'*��ggg3�-�- �F�jU���M�P��W1�U�S[�Q&�)#�O[����͛��y�� �x�W���I,�!Q��.:
��0#a�'1�t).��sQ��Y�m.��O1Gm���uq<��v�q��K��\/�Q)x�7�U��1�z/8��F�A�MhD*H$�C�N����!�9)׈�.��!��`�!.��ӛ!�6�=.�t�eƫ��߿R<#OI[�^:��n=�<P�Bf���^7@O�pW���O���:v�ۻL;�0yyi�-�U���n����Q�|��U�l�d� Q6��2��Z����l<����V=vv�-���9����W���c��l��99��Wq	+��M�KD A�����?vB��'���g����-M6����_�߸ZN �\�|�
Z}���ڇS����i���K���,;Q��m��G_[�]��Jr4�Y�6ÙѶ/�Q�9A-|CF �`�v�>{�8V���qЉ�J �S���n�h��ɒ�/�tp�*O듐��II��@�_��`c�aM�w��p1bP=>P�݆�VV�hgٶ��.��G�dƛ;��n^���5�4�(	6�C%�)�Cw��� �"�U:�C�֡��R�,2@,Dq2H�>���	�ֵ����|�{V<�����?�P�k��]����ό�ĈJj��9A4kB#�~�U����Ҿ��@Ȩz����m���,�k��\���n_;ͭ<�Y����*���� ��M|��cha��7B!�{M>^�w�E�}�`�dp��$ CDU���Z�c3BǏ�{>4�uE�^�ﾠ�מnk�����e�}A��~��q�T��ݤh��
���		CC��|4��GPnG�<`=���Pl�_d� .l3��V�x �֩SĮ��<lJ����m[����se��V>���ϟ?3��]]z���UV������۵�\�
�Z�&d6�����p���U��x���p����!�51?�al��*�a=C_��a76Bw�[�
��Ĉ[K�9�h�H����㶹������:�{*�~��y��Tְ}�˨qfx�:�-O��S:�E���WX����b� ��5��	7�t2������K����e8nS�`3��7�^�?z��wj�؏�r��>�Y���m�S�&����(���l�ʂaCm�a���;1��4.nH��ǧE5�r��^�v�ᙾ�=������g�Bj}(M��;����/����)�Kg��u�d��}@�����e���C��G/����婥�ú.��vo�U�$H+U���oT��/22��%���Cݼk�*4��zs2�?w�Ff�W����c�h\�4tuOO�x8z<��U]�L/Cw�d����ݪjv�55GtM���`�{������LpD�nGy�beQ0Кg:��*����ط߲.$)==H�@g�0D/�˽-�����}�F cO���tn�����0S��X_{�Z��p��f�N�2�{�La�3��5ڤ<�/y���(���R�*���=0�Uh�>z�� �>��Eb�N���
��N�x|MS�y�Y۵ڳkm�
(���ԕ�,*����U��+�<���T�κڦx���_�^W���2e���l0�.�~�N��/��s�<��qip q��t@@ z���o��ͽVaO	��u�?��.5�t���S�Ջx�n�;.��)++kٛ���<�0ZҠ@���[Ẍ́���#z��
��	��3]Ch�Ӌ���s]�/mx'G/��ItC�.ٍ��4#]]]�f�8�v^7G�-�����|��˨-��w�5��N�g�3��ë_2^>N�-dz�<����[=V�d$����;tm��l` �2�^�����w���6��;i���z;���ӝ��A����,���T� Ak9���4�<�+���ѳ)���97�4}�[������>��Q
��|���,��5���-�q��������,/�}��|\!���cgߑ���uv�>t7(��B��XE�z�l��|�L�]^�W����u���t�T�Ա��M'����!ڂ}�*�Ti\�^s�v^��7�)�+���g~j�a�D�R����K�?�s�ɺ��	�#�Ú�[~]�R<�a\�E5[P����]ގE��E�ޅ������vEZS��Hk��؛L��?�����'�G?�����_��}�Y'p�:�w�3�\4F¬O��$ H'^.��.;�#�?�ӌ��D�C;W���km0��6���a���7%��޾�˚�~~�#St;8z��&$!3�#���d�c����Aŵ�
�Ϲ�0���*�f�Z�Ɖ\���`���;��[��������?�Wƹ�w8��hT��������}�5
�>=����]�&A�u��~c����nU?.�������y��{� 9�+������#������k�:U�~�]����_<�����Q�6,�D|)�D��؜d@�zw�K�)��'�o�3��s�&k hFG�('�^�t��R�@���I`��n�p����A��9g���y�rl���伤�ï���R�<[Le�촵p�E���Ѯ|��[t��c�/n=~��?����'�o�ӥ[�+���7ٰi�P�L2*e�Ts�[ý�Z<{��>��<�|[�
��8硱�`)��72�?��!V��b7;4�u���?�1��ѿ�&Dx��z)�
c���d`_��3-.������2��������{�{Rr��ߔpSj��~N����I))k79����r���:/?�%�e؝�@�$�&�ᇘm5Ԓ���E���{+�}���$��-󺾼8'~�ȥ��ۿ���;6m5�*ċ9%湻�_��y��Ɲ��������'��2��b<��}~���|����5ka��@�s��,wA#�nw*�zi�n!���lI�w0��?./6�ط���m2�6)�8��̾��Ջ�+t�4�;��ˬ��aP`2�n�
�������Z��V'�P���TY�l��ٻ�5ϳ
.'�A{�}������Wq!�m�_U�lZ��ք<���<44to��'6_x���$����:	�#s�Ck~��鸻��yYE��Ov�kK�i�����ǽA�~�.��0�|��l�G	$`,m�	љ����|���y˙KT�W��l-:�!a�YDVet.�"��B�#��{��O�-~um��ws#��uu��̳9�����^��IHAW|x�`�R��S=��*���r�S�+{�P�����F�$��އ����Zf�p}�GË�f�~�lo1��;��8%e�����|&	��-�Hb�zJ8��4S�a��}ո�z���3�Q��k48M�鮈�m��9��/���~�zh��F�9K�(�[n�m75w�4��N�S��1��?7?o�qo���w	W�+g��=`@±h(ۘ�y-\ESc��)��4�jp�mO���W����p��	E'Z�o���-��Ou�&�A���P�ӛQ����g�)>�v���!��^�����g�������@l��#AD��3�N�d���ߤ�b ��]�ۉF�G���<��o�W��<�077W�c�� b���(��]Y�6�oA�g�Y���6H�?T�>�Y��>�?��+�ESSS�����~V�
�ptt�`T�\�깢�kw�:���1%�HK��V8�;@����Ƽ�<n~ni٠ZT
"��$�zQ����������k4p�����N���w�~nFi4�揗Ē�#����D�����ǈ�k��>��U\���TP��V�#�n��}�;�����{@/iim|��>Z!0�����X-z�x�-3H���N�D�y���q���fߣś������)����!	������A����(��k��Q̈́��N�ԝ�]|	3���` Xj\i��H#3]�	 �cz�.���7�v��B��mv^�_���$u'z��U���ݻK($��k�37�	�xw�Wa���E���E�ddd�<���͵RS�O���BA':�r"N��@BO�O�~��\��v1
"ख���R����q����A���ٺ̃���W��Ӈ0Y	��˚Yv���e|6k�2֎Us�<�ca�dN)p���Ɨ��Y�mG(�s����n����Y:�\���κ�I�/I5'�3��e�#��Ц��� j.�A�dO����{Q`tt���G�6�E�X���e��M[U�����������h�(�aJ���0Ҧ�TFi���ě�QV���1���R�ROCK�w��ܽ�>���>�w�}��u�3^�s��\�2�ˋ\���-�ca��(���򞈪�4=���=T�/mQ �L c��p����_�Ekr3`qk���>{����b��ˇN��g~�ipLĻ�T��e�V7`C!�F������,FW�6���Jqߌ�ˌ��I�ɳ�t���WڲHY� ��x�7���)������!,tV��{�_�������}����N�fn�試��l���y2��a�C���BCw���XvZ��g����l�0V��
��J�<��lK���>�J���`f�&e�KK���H����]U}:��	kB�I��փ��מ�����!l��������KJ��eN0��Q+��A�!���X?o���=�޺�^{;�7�.��o#$9�F{��2"~N
hk����JJ$2�� vg�=���+ PRR68�9�1z�\�2�y\������n�;�?5X��%ڶ�W�f�/+��e��b�]��2u�Y�Ŧ,ZK��D���dI�7�6l�P�sp
0Wn�+(4�&��WCM�+��!o�+���+�%jQ��h�x2˾���������+^���B�{�(����W�T����HhS��漟���3�'���+
�������m�#�*��̸�	�.�z�T�q喰� ����1�N��L�K���1��c՗�.�Z?��K浫�P �*�Ū�����{+p���	&6_�k�<�� ���eљ�t�...64^Ŗtfj����1�"ZXUUU3%/����Գ�Z+�k
|^t��$�����v�����'�繑�z�����Ol��2=X�^���*����0����@WO�ċ�c ,^csb� ���o
s��9Ͻ�=���4+:�O����y��s��D�������LrmaK�wû%u�5|�����=\���J�u~",0��������l�:�nѭ���S���t]!�����������
t����R��զ�gh��������C1�W}�)V-Fͥ��q@�e�
t@�j��=Vo�١��L�\E��/ɪ˭��}7�OC��{vd�cCֺ�2淸��Wm\�,� Zo�5@:���Y�|������� �˞T���{e��ʋ���v�M���4&U*7*)<���2!�ϵ������pN��Du]��r>qlI=,K�N�Ǽ�� �ڴ�D���`!˷Joj�YL���I��������5�^��x�4�+�'��n 舐��)8��}3���0���UT�^`-�$
�zUṨ�F�Yv��j�dp��c�G�*�M���!�k����Ooڹ��L���\]�ڕc{f1i<4Ћ�z���U���7���պ���>=��Ww@�٫- o�.��W!�ɀ`eJ��; �WL�������\�D�ڱ[W�'��.e���VK�v�:?�^�ݹ����M��?VvE@�!�͆<�GG�V�廱;7B!�$ھ ��ڵG��}ʓi)�C��j7[��<��QW�h�tt�.��ꧣ�Ԏ��Gk�S��l�>e^�@�'�q�YA�i�|���\�k���A�����N��9��֊W,ql�ZV0U�4բ0R������-w��IFV����B�K��֘�"��N��2U���8яB�ߖ�c��Z�� ���߭(u9���<ܗs��o	���S�+�K�L^Q�����Ou���8Ƀ�T��l+&�^�r�ξ;�۶%��x�0����F?��c-38�#>���B]ѱnᜇ3n633;?䚸Ե����JrSik�����E��!��J{�g��\��
��p�I���>����֏}���6�4pDE�>_;���":���??�}�Q:��y�ne���`oח�f; ��Qv[�����;��� mٶ	Ǟ�?�^��m�j���@uhNN��bIk�t�\5�G�/C��]e��.rC[��Է ���:::�{�끼;7��+K�F߸�^��˄��edf�v������Æ���&+�/>���./ebW=�c_S�����/�щ������O��W$$;� (�ߡ�&}��]գg?���9�t�+���m޷�x��iͅ�����" 
�+]�ќ%or��?�'q�kȶst$s�%�&ԧ��Oo��Z�����1�	`���9���������0uk� �X�l7�)�y��ȝ��g�`��&nވ��d⽞��p��=� ?��/�����f�VH7"�×<1���9��cO�D�ȯZk�`G9K�f�ފ[m�L�A�غߓ�ԝpJ/;��p�<]2����y'�y��ܐ�_��-�����+�� ��]�d�{���і���\m-�3���a�]LFD�6�.oۘ��"��3`p��2�E�w��[q�ԗ���X�m,3CQ�$A�-7�;��b]����y��Ú�`
~'O.�LbZf����'��N��`j}��.$$�~���OLUm}�p�cݩ�3�6�ᑑ-wo������7���
�y�YZW�����	�gw�T<�����7�-�`ۚ
��X�%��;���͢i������P����s�	qϚ��H�b�S�XE(�Y��+~U�^���To��Z��
U��B�\Vw�����B�Y�-Y��2&!��b��}���,�F�iۯ�M���f��e��e���l!�?�S���-�����lM�u��n�����h���U�둜@''�]��q��).�:Vw���S� r�{��7�:��n-XS����y^�g�5��~�k�_}}��ͲOP��o�s{�B,����=�
{\X��U�;F���b���
����B��d�,�!ZK�<����7R���� kƇ��Yv��`Ӂ��Fj�H�z(�8�K)�ו�:0-(�����>ݪ&ߤ�VMs!��%cD�5u�q��y�/�X�������Z乮��>*y���������..^)��=y�^�]m�'X�g�	�"����T���ܼ��s������#i�� ǗCL|�eO��eB�[@[��s���$7Wf��v�R)���[�M����ڶ��ȃ��mmmIakW���?�5g>��T=$x������O����8G�my���c��6�Zf>����xGXD����lO	�5)ls	Y^	�y$��˳�J:�������s�#*"[	AknM�_Ӳ+���v�o��L�q���{{Ӛ3φ�{?�ہW�)�l*�U"Dw-h�Y'F���)Wo��!yâV9�����tǵux��RPP���*��j�N�}:�������c}�N���cpA���y�!�*ǩ1ø�{Grƶ'w['$>ܤ�_���S��H����jJ����RX$��{��d�N�N�h���o��h<5�߄�r�)n +9_�J�=��\���Nyr��M�4Um>���ڶ�D�I�2o |���Ƒgu�c^�[�'l��,�:;Wx�pn����d�o/. UIII�u��2a���w����_�&�SD%�*c�}�]���7-BCC�=��t��/�]~V�جވ1���s�V��3�4ˏI6;,�a!��ĩ�WEJ�L_)�wGPk���d_c.���<6Ff��y�n^���ј3�ڀB��Q���QP�Mu�ᝍ�ԃ�����z#k)�"����kMx���=R��u]�8U/g~�7�V/ޘC\4���Å�A�mξ�.����clX^Q��������<�U���w ��C�^�*��!�r
���U����������h;5>xʹ{x$������Ҕ{��Z�TY�3_i(썡�Q����$F��~�N�{������;��Rs�=��p�����U�L�9^��os#5�͞%J���T�,n�qP]�80�Q�����Z�b�����J�_�Rv���ٌ��Z����L[C�w�n@O�������J]�~�	���	�@W�
+ɼ��ϝ�,�-�xB}�[�����Ot��@Pt����o? ��?_Ha�^�p~ǣG���}4[@�R�7���X�y�w��R��c�4�����SA]���,I�_np��ep�O#vﴰ��h���t���Ã�j �m
#��;����Q<�=���衁��
������]~�`d%���nK�m���j�nv�/�6�-���fܷV�]��30cU0�%Ď��JCb��7}�����6G����']JE@��S�ِ��Z�n螯���ڎ���^;G	���r���V�|=��v���w�LG�.�C]%v_�?LMM?{/�F�b�z���Zwߍ2�D�(��B%-��[��]i6#L�,����κ�b�IO���	��8*����W�����RiE�q�W����8������2Nd]dV��
sJ���G$]%�@���Ip�������Xݥ�H�ݪ������k�l,��c�pH�����19�g��MR�o�u�����Ԟ�6,
�h�ehw������/	�z �����TjEL��y�6M���,��i�o�%3�,2��+�'�ƴ��r��(�R���]l)�r6O���7Qr���3x��H�������W�9��� �n���Tƛ�]ŹϬm˲�ʸL�2yz	@f��{����ULrF\ܫQ$�@HX�lEJ=����m0��c͒�n�.���D�N�+4IL�f�2`��=naţ�2�t=��mi� ��cog}r��ޭ<0��hQ����v�(���²uw_�A��$����PEJ,RJ237������L"ڑ?ӕc���=s�;b�]7������^���\�����}��7����^^��|A=%�/����sK��&|Fԥx$�_>�0���{����^)�����R����ݕs�->ĪM�����(kᤤS���^�/����:��������ǾNN}�� �7��/6�����,�zG���K^����M��� �N�fy����R��?4V�
�:�' �P�jw�>�;w"����Hׯ_������;W�k�N��<s����q_�40^PX����RMM��"��!��?����e>X[P�k*����H:�������r�x�80U:h�Cy�~}���hA����j�y�Npy����uy��:D8���Hi�8���PƝ?Y]x}��ݙ���:�DGUd׮� L�݆p������E|�zfƜsب�ϩ"����HP��W�¿�Ku֝������W��8Q7��*O�B�%b�A%��'H�EP<|�WK/���S�7��@���&�Z�����i�N#��y����_Qч�y�z��'Aa�kP�9���6,��_��?��c�Wы\f���'ڢt&��!��K�?�\�&���*��<0z��y����s�O�N�њ	B0�}�� f��?�+�G,s�ul���ȋ��-Z���1�5U��	��51Q&���8&���`����cΚ�(���Ù�zo�:0��}EA�� �� �0��oN�S��r�*��8��?���M\L�׿�����OLϘ��Luq|�H7D̂h;��E
���M�X�v��'�G� ������~f�Z.P�{��Q#���ΐ�#[��R���RQ���0����� r7����b�_�m-NX?���kz+�S15�{*��)[1�I�����5 ���#JʘnX�FXSȒ�������
���O�-�ey �$�N 4d"�4���=h�Z�L�6u����OA^��м�^]}����W�T���\x�j���j���eR~�GAJ�����!��4(ns�B��V�aI�*��!��5�?/�[=S�(�%����a�_��	�����<��Dv�a�#]p&���bՄ	���s9��I>@���w��6���"W/�9X�)X_EP!��e��\�d�.!�7��)y��d�vb5`��G^�CA3C�]V � ���ʰ	���.�"��~�b��z���	���4����2��ԇ�;0���{Gy#��	̏��1��ﹸY��l�k@4�o����? 4�$f3�HX�>�B,j��E�ט�q�0���A	�ډ���>�6>}�4�ſ|����d��bB�D�o:~R��C~�z����й"a`yso�ٔ�� od��ػt�w�R�q�?_k�t�J�b� �Iy,QP�td譾L~Mu��bblt��0�I�e(�������l�O��f�85_E�r��ޞ\��ĉ�摮�5��P�n��z�M�#��s��<n���97��05n� 5a���~�`��w���J,4�*��ݲ����ӱ�<l�T��nc�����jZb>lx���1�!�y���U��Fh���8�R0~������Ǉ��<�F*Um}�m�9�u������zŧ?�"*R�`l5D�]���reK�wkD��k�������0+a 
�ڋ�k��Nv�!,���ss�*1݂���w����4���m�����f��������y(��F:���7��o/�s��h ��Ađ����~,2E�����6��[�^���{��JƑa��~"ޜ�'a|�u�����Vp"u���Ȩ�<��1�8FVX�F�X[���O+�.b���rmccc�h���f��$|�������&�o��tWl��K�&X����9��L7��1?��7��%1��0|���m�`�(�w0V���b�� E;��-��(9v}�b����\j��Kh�zb����
�d,J�=��߂�S�D�'&& ֚�Q��!(�'����/��=�)P�|�(˰~~����=|8s�f���A�{c@��庤��Z.h�uj��ege!��\4�i��<���b��9�r1J����nT��)�6\�..i]}	�R;���h4P�`��f���є�SCV�ߟS0�6�M��?N��;Qa�NlZ+]��1;ݘ��I�b�'9�X6Υ Z�)��N��vL=��[,��߭R�N�tc�"�-c�)��F휎t��NI%��R�ً�$��l�T�
�ܝ��y���[�<X�I��V~�&P�b�����Ƴ\"�������h�$��3~wqW��z�9�v��W��Aߗ=h��+ƥd���ne���N�>��!}��(���'U�������~�J��a�R�mhe%��ܼ�����^+R�)Q��G�o H˟,���ϭ���b��mE�
 �)Ve����� ��(2�Xw%.�O򧶲r1F��jZZb��`��:^+Bw�t)f��9ᣪ��5�3f�iM�n�.àˆޖ���E.�9e�:Q��٠����Q���}|<����TGG��Z�8��^���$��jp���dn���b,�ؒ��,֮����|���掩?�a�;T���\a8^�v<(,���ړ�N������x�0��廛R�k�
�we�`5�QV"\�&֕�c�<���ľ[���Β:���[b��:,ZY L9$))	k�����Wq#+����c�L9��0����y�o���oU�"�u��Ö��Џ]����+��l  ���n²��̊ML�W�5��e�f< ��~<Gc;1܍�?(X�#���R��kjj
c1� �sr�~�=y�iWfÊUy��i��>r��=��-�m���N~�@CV�EL�X�ȭ�m���8�W�,[���R]��ޫ���^-���S=�ՐI_n�!gl�����Eߣ��y��8&�����?�j�|&+�Y�uA9w�ণ����E`1���"�Av20�z��Z��j�)J1y�L��߿���v�ݗ�<���᜵g���m�'�=P��Ӟ>�.p�^��3"�KzwUʰ��x��;��/��^�,�\НD��n�,�?��#�g	�9�^2�Id��O���3k��v�b�d�!�F���qj��r�5d_a�Qg���0��١� ;�\F�7oj�]�����/~{������y�ӯ�]�6�q�ki]`<#�x�>�~��cz�jo��!*�%�M��q-۴Z�
ș;ץ���&F�4<4+��`�PZ�������/����F ��������g�����ʷ���.~~������`�Iʍ@F��_����fd�qI�d��Xe���h�TA�ߋ�_�~=��e�_�t5埖�*�JP
6:�=[�~����iB` �7"0�Ќ���}��i"��ܚ=j!x+�
]�����<[Vc߹3��c��C_���:��yoit{ɭ��"�0�gwl�x�ȅ�c-6A�� n�o�oy9�Y���3��^�P�o�"�C_P����v����!����O��,�hM�0~,>v#*���c�B<�D'��1�.�����ϴ��]���K�V��Fې��:�"�Ju��ugg�Y��=�7S{M[��a��oMk2DEiRp��<��  P��(f�����og���׎6{���y��q��?W7F�<�E[/#z���2��%�f�Ɇ,{���oZ��:�Suzf��x<d�f�Q��E��X3��S{b>�ݻ�y�&UdF�رcM��N� �`R��d,��:�}ϡ����˪H�C@!��L�d���ܼ��JZ�X<��.ݖt��A>�^ųW0�����a���/�	�w���|��F~d�Z@iD@�0�d�#�����޵0h�����L����*�N�=���@6��~����P�Yn(;k�j���y��-�`q�>=�y|��7����	t�6��A�rr:t��������w-��b�O�3	�h����oh�h��ׅ $$��uUppyO;`�^eee��7��Yi�x�o�j�g}DX��L�#��y/yF��T�h��G����W�o�t8�q�܃߿�R���������m#��P_�$��e)�����ME�����h2����u xea����ٶ��k|���\��7���J!��ώ����FM�f���I1+�zb���1�����>l,u��b	A���'j���8��UUE��^����i���AhLSw�"%T0�R�1��Bg�:��cm��/�����B��&�<+͙�6�,`)�b��1����u�f�dԖnp<ý��)�|y/� ~��j:�J�^�/..*����#��r_E+80u�˗�ޗ��5.�ڻ3Z3�egjA8f�T���}��0�Ɔ�������B�W*b�e����=�1���U@x˩�YN�d�˫���w�������Eԃ�1>�r5?�v�W��#��%��!Nl����D����j��l�)|xvv���3݉���ҿ<��>t������w�Z�q�I�aj5Þ���^u���z!�*/?��$��udg�Nc@c�E�yE�S�����ôfU:F�&#r۫�C��Ե������W<1a#��L�X,��=�&`yf�s!�ڇ�O.AM']�U%��e>��
��| *������J�5c
��g/�!��#�V�_�ϝ�:Q��zv�z��=J���B��m���R.vv+&���~4�%K��*�^Z�����cQ0���W>#=K���7�@��u��pn�)B�$Fݿ����EogXb7*�+ܸ"�'�,6P,V���L����L�b=�g�t|Ɖ�ع�\Cb�M�`�Yզ�j����//�27��
���Ç��l�S�yb��՘��vX�P@��&<�lF�kii)��wW&�c�{a�S-
R������Gs6�K� �1"
Q8+D�N����u���-�pSt�/��O�;�K�'Ac�|���ͩ��� �G�~~�ky%�ǉB %���|;�� �u�X� ^a�dy����(o��2-����d�%��'��PYlڞ�ϪV�׺"��ɽJ>�ة1�4�Gy�����<Z�/fB(cW�P�[ɸ�����{�>�v��5�}�/yg���&�:������A�w����;<���&��m�-��J��y��u��!]�K`LL��U�Gȿ�J���ى4,���B��`���ڋ��k<\ ��R"-BOeEM�5����P���n�ϟ�i�lhdDR�gO��N�h`;�q�b	��?b<���ג6_�Bp����!�xu"��o/U�/��Ķ/�O���+#��8Q~��o0&�6�i[�g<��2�oV�1�PF���}�jJ1h���\�VP�K�|�D<*���G�C�F�tP��>��o�&|S�Z�ju���'^�!��Tn�a��h�U�����:a��ֳ3��!�삯\�H��[�3���� #�d�;���\����l���xn��ñ"�!�IXsda�a���4f����=z�X1��0򖼽�������<7��b0�g��[��"<� ���I�iz���Cx_5����FT{a ��~hH|�n�Qx���ǡ΀�cQ�gď^��ޕd��#G�z�n�
�8�/&�C̚�x�}�7�[�PA ��MB3U��?|�-
=I)+���6�E�<%�E�0��vnVA��9�c��-����nzX��M֏C3%���f��gp�WQ���>�vݺ������~�X��4��۷y���yT�E�שN j����1�MKe��$gdlBר�����r��t7p�Dg4V+���@��?����;�3V�Z �"}$N�REN����I��Dg�U�^�o;O��8Y��'���ϸ0<{N��.���[����*��z9,^���LZ�|��{`"<R@vA�I�i�t�<Rm�q��L0�f6�3c!@R������t_��u���{�Qu�bͪ]eY:�iх������/�Y (�cOp���7+�@c!����� ���U��0ar�=��q w���$����p�d,U���ɻ� �+_����9�GM&��F:�m9��f����Д���נ@iX��R�e_�+ۡ�1aHw�9���%n��Z۶�;ך2	�E�� (�mw�U�y�b��?,�@�����W�n���O��X�g�&�-�}�ɣ�勮4|��4W�輦W�uX��e�x��B�<�p�+�R���S������Џ*�:VFY�Ô�5�A�݆�J��]� �ӘGm��c;���|� ��ݿh���Wg��A � >q�!����=�F�s���s����p-9��_@'� �B��x���q���"U��n�w�YUzW�Ȗ(�f&� ��>�dN���n.�	��؎��ԟ�χ�a����U���Qj�;�b�ڵ�����i� MDkB��f�o�%Wg"��uF�Jc5�b�����wkaZ���wٳ�:3�p�&�L�R�?홟T�d
�����hpE�𿙪7�v�g���
��	Oq�g�@��E}I�����=5����m�{��7ҥ 
xjC`���sx�΁c�z:���^Q�)���iU=�g�%�j�?)w\]�����2w�my�?9Z�z�L�������;���_@?I�����\bԞ�,??���/����|�4�fwc����ϬƐ�w�чLt3�.���#�#"�w��P��ϗ��	�P��>��u�UW}�	R
;"�6齌�C��蹋��`��й���]w#�?��IP*6lSF��x^�1`��;�R�G�.}�kY>x��ھ��披x�P���t@F�>��������9�	O�+K7�|{q��,����k�jLK�n��fD�:�G�����$�����ʰ�K'R4�}]�wA��WO>Q���O[�M���
�g ׽�� J3�!n���
>X��/��=�g��]��%�Y�!��J���|��g��2?���Xu�y*{���9�茩��T��1�:�ԪT�h���܊���K5�!(�y�YtT�iz(���2�x��!Q?��M����vle@�^���71�,>�Ez�[¹x��/�_������e�$�y�I�w�lN-�������.Eة�z,]~6#�L<(��sr�39������+��E�3��'+��iq� v�,��#//�eg�\�з:V���%�+�c6�[E��N`��OjcMv��� pB~�X����93�-^�i��	���?��O��7V�6��'�D��3U�2{ىW�5 V2�u�v� �&".Y ĭ�o�g��!}�h�= u�Żu�iM�`��6%;�P��:剮����K�F����E�w�*����%�Psz5�o������n��Bt=�)�PZQ���u��~#O�B��"�T�50xn�yu�葅Qh����}����Ɍc�)����؄���;^-�0N�,aW�J�C'D�Ā@^�~]�������2l�BTk�g��pyT��8M ����8	�$����՜����le<�be�=�j�u�W7��L�\��t�r�٩ߙ���5��Ua[7!�"��a"�x���_��`D��jK�����7h��j���"����]�r��0�<[�&͗�uG��>���b�Q��w�H��`�@9�"!:S�}�&��oP\��k)���ո���h ,og��R���:��U0�ہ��}�r�O�Dg,hG������4��U��~�~[:ǹY��և�p^�Ζ�~?J�7#�-��ك^ŭl�)#v�v���[A<������PsX�`L��7<u�9tB��А���k1R�����[�o{��;���r1^��$�&��(��|���&*�ڣR�T�B���l@X�n�p���m�sͷ������L�ͻ�&�.�l3���\���U-p�����'+����Z�n�����P[�S�"_ӊ
��K_��n�0꼀8i�#n�KL��Q
�J������ql)�B����A@1�?�(�1��n���)�y)Q�~O�������[�i����أ�uv����En&M�e*�v�*	��'�w�~!��_��x��ƍ�B�Z�q'�76l�mXOZǩ�m"�?��L'k� �d#��C#ܵ�3Hڵ5�>�*2Ԅ[]@�ݾ�4Uq挿�Y��;] ����'C�9�9�*�rvv��wNLu�����f3�̭c���B�/���ek���Wr�Gg;�ʠ��]J:c���^���t�u������`%8�g��d\96���)[$'S2�>��:���-n(p��Q�܀pO��9� ����0S"���Ѓx��A4Y���G���Stjx�T2�x��HԔ���æ� ���&�;XM^����u�s�~��R��G�<�8#��t���2�n�?��e������ә�%��/X
FY����������U��LE�рD�$��r�ܣG/�ڄZ,�,?$�t�]�Yc�ǹ�|5-�.D�/�m�8ỢL��\[��I<�����:��Z�:9�f��_w��R�K�yT�΁���� �oDE	/�g��(Ɠ��sW���[�1�V/[�/��� ���5�!V�-Sų�V���$9G�����ƿ��-��P�R:���V����n2i8�	��o��5��:���gV��e����n�߄0�y��z�ҩ���/� �r]Z���`أ���q��8b|���A��?�&z�t�ǚG�J�Ǌ�x���
��K
ho�"�G�Bd�z�:��P����L��>�!1;&1������Đaö���/g�IN�ϱ��Q�n�fƕ}�B����K��Ua\����N ���`W�W��Ҋ*�{�����uC�OLR��q�\�J�[I/�h����\r\���SoV0h��4զZ�R"�#�t���(q1�J���#!hV�K�I��į�; 3p/�
���� �g�����n޼YV[2�����C&������(nx}u�\S��%��ps���C�NC$m��/�����dz&#kEGPg�n�)��g_v���!�,�+�A���x�/� ��%�"�燡���!E��4�A��)�Ω�T^8��=X*ϕsh�sm�bF�w5���Z���K�b]A��H�mq��Y!+M3[JV6��X���=�O;
��hK�$kS���1;�ם�]拧%�"N�m�%F_�N��_�`�7�0ݪ���SQ���J���׀��Rt:�����K�	yw�����:t�Sg,�A��H���B�~z7�<�xeV\sS����;�4��e6ϔ ]�s�ao\[$ȟ&�a�����:���3�y�0�tp�Z��*�`M��x?hX��hn:�������v�L�R�/�=H�1�
~��]@����J��]�Do
x�����5)f�}ه.-0h���	�Cy�ʒiOCnJt^�v���>hg�����â}dwF��WcJ��)d�8��UGG�%^�o�k��*�pO������9&F�"z��k
�� 5������ �^~�-s�C777��t��m��x��X��X��\�e~���`��������%�����a�J04G��N�C��p��O����}���L�,E৾c�A�C����/�f��U���������ڂ�$�vt���W�����d�J|�~iU���|ML'_�`�}M��b�I�1Kw\�z+S����G�H0��VJ�skD������]�2��ߢ�K��L��y�ٻ}� p�ܹ���]z*�����0̽�%1�xT��R�13j�ۗ�n�x�B����###�5uu�
�"o�a��ػ����zLK�q��5Q}r��JUQ�i2�+n�-�U���O���߃^xB_Ҍ������/�!�4����������7�A*��n�$
�]]@QǇE^0��+7��{��铘ur��U*2���gL����R"�;���q ����2�
�80DU��.��ث� �����0�-	R�� �X��ľA��͇[� ʣ���;Q}�0�>'��P��x_�[Ogp�3�9��եE�1�S-g:B0d��� =1��l�*	`�E��Ӂ�=�k$qr/,�M��C_`��C�8��??b��k�l�?���w��;��M��j �T<Nr��I��T�5�U%�{5{`��������@֢�.���p̊E\ ����E�H{�=~�@�T��I;��n��IsG��+�M��b�-���֯_���19���[^�r>�ȗ���W�=�k��Z�����θ>�C��nܼI�PM���4+,��U:#�$�.�Ɍ�ME��GO1#N1W��LLa�K���N�/��2�������Sbv4�4;*R��Kf�VΥt uL�Qn}�)�fX��!�1ӷ���Sr[�����i��4d�3��<eB�o
4G�8���_�����ԩ�}�$ʹ(��y����P���3�¼�m�>���ӿ
#��Lݳ�!W����Dm邦@�5}�7߇aTV7��LP.b�i��y��1�%K��c��y��)���5��M--c�N�_�����:�%���ޑZ�
��Z	��v�aRYx����<�����e}���sQx>�ʒ�<ȫ��l��K }���G�厜<��ɬ��O���QV��çO��W������k�2�:R�j����?��X���	8��/��b�$������(���[0��:񐷒2��|dh�m � �$T/��N�[Z��GJF&B��!r$�^��Yd���_���R�۰��n��ӻ�¦���`���g[�����p�����Ƞ�:��8Fe|9U>z��\���3r�;>:a��=��ҢU����x��{��1uoV�j�G$��薞(�LZG����ܑ�0Y6��w�g	np6���H����B�*�|��bǏ�P,ۖe��	�m[���ڢ.0�%R�#ԕ\����X�,h���nL�Q��O�_��BR�r�T�����(��7�V鞱|f���s��1,��L�s2_��l~UTME5�)^]�|�F�i�1SK�5���?~o[Fbǀ���<'w��ܐy��}}�2X�Zf�Ut�?Q�؞���6�X>h�e����Y�U0\�+ǥ�О=�nxz�q�����ϋ��riU��t��W�߿O~!�&r�-pp$�Z�ٙ?���́M7lFW�*�U������}z�5B�Ozņ؂;ӡ��,٭=���z��FbҚ�G��њ3����[�G���|�2[�^�[���Bg���}��uX �v�?���"����cd��*�Z�UT�V� Q;$'��.�ss�-И��tkt��Sf9�moo�+ ,]�8��gV:��elX L�D��-q|N��~7;��.�j�#`{W��u4y�鼁@3��xز����ᦎ�o,��tf�G��Oq��/�^�����(6s�Xf���d����S^�3�ܹs�_�û\Yn''�(�LP�1�u�5m��'�����}hŝ�7ݧ�ҊGo��ʹ�=���n[�d�{�����1=3��&:Tk�{R����\���a�,��c�&q��T��M\�5:3=y�<;��[�
%/G�@d軍�����O�I�P���>�[���� �<O7��mZ����O���s��'�[�ɲ�G����4����JϊQ�U�0�L��>�����̅@��n�@U�^�m`���U��9�[6�ɳZz� �._��N��� ���lW��.�����e�$�D<���scoM�����;k�������{wj}��^P{z�(6f���4��E�ar:����'F~E��|��s̘D�6^(cQ���Ύ�!,�K |�
�s<�.;1���qQi{���T������8�M���9��Vv�������n	V�"��^��|i��X��V�����V����kv)Z��[-L49OM��9{��	й�����=�>��59�>=��}2K�^�c�����13)$���5t���]R��3/�{��un���1�g��&<���g��r7E��,hbz����vr���J�U��+�b����)HS�|���5�<D������e@D�\�^pb�������㷝��~h��q2a�3���b�A��vE@�Sh(S�O�}}��z�M����1`���V��T�f�W]����S,�ԚS��hy.9�#:��h�����Q����jɒ%�6�>$ٜ��B�Ȅ@v����g��VC����<�7ߢ��mn�#0�>�_�����S���p,���^f�k�KR���urkr+?&�=�J�ˉw��&��Wt@%���#�y���l��|�@�y���H�MD6����1Q`�?���_ng:�d��'o�ƪ��J�,n�?�@d.�t>�;O zŭmQ��¬ث�b~��h�E�k����;xC@��D�j��d� }ƫ�n2{Q
�����r��[`^����%���/u�m�շ�NU���K%������<�+����t���݆��Gq�1�"���q�h��%�}���j~��ٌ�q�~ے���_'J��X�������|?�a��y�G�sm��\Hr�B,W�=�~Y���?k���/+���+�Z��;��p�}|����Sm%f��h-�e
73�ի��ܥ���MS˷������aA�M_��^���^�uA�qv &�J�3ܿ��b���Pm����<Jn�e�8Vl�]�wt��#�	Yn���<M��4�x�'O\�ד�#�~�mF�[��(�
��c��&��fUP�8v�[DHgk�m�C�4�1?=�s�<zh�{�m۶):>v�s�PȰ ��0c�iO)W��"z}���u�K^ ��̈�|��w�h�|��T.������Oڥ6��3��.쁧�aR��4{���ML�;�y�S�}��P!��_m?`&����ں���D�]@�X��9QԼ����+:��s��ӑ���͒�����f��v}����S��ǳ*c8U�B���ό�zN�>ǟ��!�t)�\X���o���m��M��9�_��h��>�8/v*\Qc���m���shc�]�p����^�s���(�tg�O����5J�&�E�C��ޛD�9<�[E�J4��Ȩ�j��lTtj�[�����c��@��+�+�|RG�������-���Ұ4��h�3��X��8���X_���f�}�op~�^�ٵe}�N�OF+8���
�?�R��jS��ƏtF�FI���}i���7�G%u����qulɜL�yם�GFu�Z9���x8V��t���>�j@�ٞ={�{��	7��q�+�,�3����ޅ"y��E�W�0�D���;�yIX,Lz�?=1w���]%�(��[]4�'k5���w(���� �q%F��z�~X���F�,�n��s&:nԁw�; �	�U9��g(�T��r��˨"x;��dޤ�Ru�N<<[9��ݳ;Ɨ?�V2�+�{y�����Ё:��}ol����
��7_�>�W�oͮ���[�>��F���i��I6��s�����3b!��a�
�/_r��|���Em
[[������˼oi��خk�2���o��ͿcN���~�f����m��%�M������f-|��2�z�N����G]����>��ؙi�}/F;��:�-Ί��ˤ�}0���E��Yư�\F�w�igU��ޝ[�b�4�D|�/�RY�XՋ�/�X��>B?�gJ�k=���;�N��{��l��6�'��YX4�{o1��N�߮ڝ��ud�2���q����q������	�fff�-œ�+$+D�]��.~�7���fd�Q��MynݵA�Fyq�����ѩ{D�>�g2lj�q���k�?y�Py�׬���v5��՜yB�g�r=W��ٙ.M}+��v ���'���{2b��ѣ���D%7;�=#(�\�Lod�]��>����{���05M�b�U>�Kf�[jk�������W�E�����皴- ����2qO�g�v�ë-�ύ��$���8�Pfn����ł-�-l�����T�i��g��xq�����ǧC���|��Ԛ����XЂ�|�+����]{zE�<�O�7p������G�˗����-"�����ƒ�Љ��M�����Gj9����H�}?EL�b���o�C,,�_����j���{��)���Z�]�8e�����Z����@ɖW嗋�I^�@#;0�EJ:���N[�Ӱ��d�%_�~���6B�����U�"��L/�Mr��Mc�������=JYi���,���������G�\����.��͍g��g&��|e�TS���bw��q��+�+#�� m�� ���@�oA}�_���Q�W�NŰ��j�?�����+9��_4�N���S`QZ�������~NN�U���@_cc�f�2-�c�X��U�L�Kss�lm�Um�K�ֹSjta]~��w���s�-V�L��F�����[�˂�`�:������{�	D�c�F�U��u�$V''���ޒXR���l�P�h�����:�e������1Ji�i[�}� j��J �K��͍��������K�e�\F@'R���B��~��I��{��kE>S�����ٵ�����2k��V�6��-�V۪��W}�Q�ʋ6����QDxKR�?�$��$1c�Hi���H2F��=﹟��9�������k�u�9�<���u��}ہo'��mHaK+,�6��c���ށ?�soI�Sy�"h~c[��J�:�o6��܀�׋�V�����hj�uq�M�Î��..Z���u�y� QKͯ�
C��T(|4��R�2jQA�S�	����~��Œ��1ej����Ѷfe--�FZrnj��l`��^=���	�������-���h0�JP�L-�\;
a�=51��0���j�vg�Y�7~��`��F����f��Z���,z
�i;#�pz@��c����g�5��{�VJ0%s2iDܾ`A�;������d��%~#�zVa!R��x��
`����4^Fj/չ�����{��nڇ��&�%Y7��Q�(�*�9+�����lE�Ԓ�,�"���P�}�a���N��a�����z��}��-8��N� $�����P'6�K�&�}>�K$oټ�eF{)UGG���2�;+;w!6��*���Y~�؛��>�����4���º�L��	�d��U�E�J�����w#<�H�\�vF^������pL�ڏw�̸w0�ޢΒu���(&�<�]8�9��Yk>C}�g�KJJ��W�pb�Ha3�>p0;jԋh�;�@I���p|�%���!��.�^��z���@�2|�YkY����A����F������l�����H%�R��S�L��̟Hv ����!�çOW�_����s4�����J�N>��� �W{����[�%T"RT��[�l���g���-�:��t|>�ė��ل����z�kG}S��]�ې�$X'Wg(y��ÇK��^F<ۉq0']W���������N�� ;��u7�t0�8�2K��PW:�mԐ]u�D���\Q�Y]a���뱎��hAa�)�{+tH��	�)� ��3���Z[[5��Q�F&� Up�y�S�����=�(At��`U�6����moYlO�P(f4jQ?��W>C���ʓ/Cp~`�	��9�� ��j�@�A$������jqL�zd_S������	>G�/5��Y�!��$����Y�2�\H�\�`���blbw��2;d�R%�2Pzڗ��Z"�?b%蛿%���[�� �&$�>��ϥ��V����iΓ���Vfe��5�(�u��{��Iw��VA�ǿ�:u�+��EP?��1�q#��r�˶;�J:1�W}�/I��tA_z���G��x��Ѕ�-�M4�� 6�j��ˊ�t�g�ը��\]��"�.�c����^Uik�IN0Q�/33S�<Js>��R.e>���G
�p����
6�
A9���H��C>պك�͑"�wATHlj�$sхm~��Ϋ���~�����/e�<�v�Ub�Ha���Zu5��z�w���Zw�4����(�`7^;�:sO�%@~V��Z_��j���C��3��3�N&�l��ro�M!�����x���~��t+��|��@�&�gI��+	��!�bx��U�!�x�����TMD�PE^���鎡;lģ/�T�����vj��4��T>��v^�G�w�5��sL��~�׷ۦsr?q��{�{�E��3Px��p6!1	���h�p���x_�/�tVö�6�VߕTPTT=��L6e;T]�)���L@<!�ǬX��ONҥT��:M���~��;-�7��@G'V;p*q���'r����8�2::�x�Ȑ��X�����~�#�Q���72l)��Kn�6���g~*�� ��}��b��G~������.P��H��yx������ẩY�|5�D�=�Ũk�i?��V�0;2�'&��$��P�P��4h��(�J��5&m<�vi.c�?��߿�{�rV�3�������i�ٴ˄1,��������ؘØ�6;1���v���O�ݭzD� �\�T��\�T� �|����!��}y�jF&&&w���cA��'�����{|�ɯ���j$�+�d���96EUʹ����>�H��ͫW�..d2Y2�
}F�4�m�c��*!^��	�E��.s�/.KK[��]��MT���)�2e;�p3�:�@	�ۇ����g6v�����%Q��JuÉC�|c��{���:$���~5���9����h�HA�����զ�`��V6�$���A(���<��:��O�{82�F^��/ֿ��0$6H�fQ�7?��)�BD���$kkk?�E�,3�,}C�>��XJa���@,#��p�Ro����F��T�(�[k].,��7|���/� ���PG�_�*y�'I�~�u7`p��ia?�'�RJgz� ��d2���4��ȁy��B]���WC4�a�B{�9]�*�t)�c��$� D�`K?
�  �T�Z�8�bS�|pR�!��*�miyt��b������(oe���(`��:ʰ�ޥ����)''�ú�聇]ř!۵vuָ͌6W���.�N<���:�b��*XhWnm�9����\�V~hLØ��H^Ae˗/�Pwm8�щ�Ɵ�+w��`rw�U��1C�����
�����'j����@dk�bE��A�A��N��Q�����P(���ȩ[;yb��5�i���=[?oojn3&�n!�"@�?9("S�[��}m\����\E��7--
 J��i�WI��c�X�7�x��ʄ:��YC�M6&�qa�J�yA� ꅸsl�p[��P���R�\`oo����wp��������>H|E@-r��ʅ"���s�:�뇑p�d���Xl�;��BT�J�<�����G��)���S����(����L�g�J��ߢ�nR� �y��f?5Ԙ�O�4dP�p�����5�Dy?q}<�|�u�����b����W�9�>�I�S���0f�b���jD�����5�~����S'Nl/*D��X�����+���a1�Yk	�Pk����ا(���o�hx�QBdO���ϻ�O)yqN���3l�xw��3��ylU����&��g�1���1�޹����ݡ�J��8s��-�KpÊ��e� )婷�HFF8��.F[�"�JCP#�D�8$۠���.����V%�h���
�DW����`��$���]����!�di�����V� ��Ѧ}��S
$�u�K�� wJ�"�ZM��K���l��Oe��,�3�^�xtt"z��[�U���ǎ�&Z��l���r�H����3� N�҇_'�n L��cE�X�h�&	������� ��~]2ɗ ��}�`U�6�<�$g�Sk�IO?�J�>�Yd~n�B	{�����h@��8sb#T�*��ͥe�ۇ�1_�a�ο��� %�,��("%gM��h���X���X>�����_���e-�<cSS��ȳWd�t��� a�`�'0p�J'���wIv���Ƕ�m.��r�W6tn�D��^�
3H���-�z4m:�k�_3s�)7vp�=�(SZOO��a�]AA��ku��!�0m��+� F�1�j�>�� )CP�C��}�����xzR7����_���c�d�f�B�@�>��~�`1UH��6<���S�p����O�n'�mbon�%5МG�jD2���ai��!��R7%�jY���$d"	��BD�H���u��GNֆ�T�(���z����t1})p�jz�nʆ����tH6�l�P�� z�p �y�H��҇|��=K��ɹza��)btC���C�9{	�˳L$���Q�7w�^J�>����9d�d�V 
z+�)K}���	��J�� /�5��mȮ��vaR�������j2��<�1����c��8����6j�H?�"�-��v51�@�K�xqfMAaa�S��.�k�*<>�5�cH���及��Ď�Ϙ��dި�w���3�G^��1�Tz,<��Щ�k��J�&��t��PMlG�k�� d;���j9[Y���YZZ
�J������QW���7��,��]��.�&=�QO��B!�z6��\�1��xl�	O5�sͯH��gVVV�?��Z1Y���\} b
؄0�̼<RbD�t���,��{���?g�!�A64d�wDU�e��ww��RG~:bː��u��'!K����*�e~�` �E�N�ǳ���.ޤ#���x���p�{w���p���D���ϻ�u��4�xcRkk+w���v<�s"���i�@g##b�4b�xQ(mo��[�ͥ���T\C쑂�V\�kҝ]	J��� ?�ɟq��_�jmfW䱓A[+���x�㛞�!�ރY9�w�^���"N��������)�Q��:��!y��Ң���zh���O��1�L13c-�^9�966���-ǩSy�)K�E��6q7#炳��ҀC�2Ǔ����Ȫ��O�:zja�m��K��!�?R~D&n�ˆ������o�J�L/)�r�#�!������7�2��4[YY��%��q���!�;��+�3�y�x��A6{�N_t�:d�@a༼u���^���x���NRzv��ߵƌ���i��,��^��7!��Β}b����O����P{Di�j��g�ͦ�ih���j�6ܓ�Y�<H�-53�[+"xT��'��At�=�[
�Ό��s]��s	���u���a"�������2�I��
'N�?M:��=x ~���n�5C?�����-aK���-aK���-aK���-aK������VS�7-�/"5#}B�j�]��f�k����-�
2���*#�8U��Ob�Ÿ�m�<���3>~��9>��9޽�
�/8/w�I,�݂�	�
'N��L�_}�}]�cI���	���#6Pb��(������Hг|��F_pE�Ρ�p�F_L�34w�iQ��JN�w�'�������m���PK   �}rZ����  �  /   images/a36c4c40-5e17-4d78-b145-5ddca5d02051.png�W�[����%�0�HǨ�H�tcа!)�]JM��5i�)%����o��y�=�s����8=5b:,,,bue����@��� ��?y������m�l������S���+���������[w���������#(��������
�02�}X��t�: �W��^�Mc����*��?�\/����;�~�*[��aQ��������H�J?���S��.N��oC�ģ�~�}����Y���b�����ǭ�o��k�I�)�a����WE��q(���_2��_Zg$'�T��y1��W�V��D�xVn����K>�;�;�!��#/��GyȎ������	�KŇ��Q77�-�F���Đ�L�&RN7��Eg�-d�$��8��''���T�@ �7���B4�wwA��nt����AAr����1=W��^l�������P��� �sa��Hz��N�[�^e�wc�a4��F����k�w�a&��ڷW�\1=�H"�)��=X�W~�s�@L�r�S��������N��a�W6w�Vrw=6�s&*_Z�G����"�����1����}yyy����)�:݇��L���E푐S���Z�7-j��qڛ��5G�|�y�H��^�ٝyiS"sܖ!�H���Yc���Q��ؿ�H�H�N��J����ৎUOPJ�%��<r��֯�宭���32?ڼ!�^u�x}���T��v�˥�������j��ꋧ?|> ߐ#����onl a,��aw�������z�����z,kjj{��g)Z�'�������2G�l����]fJ"��:ɮ�C1��TT����{������'�Dd���3�t�N���ϰ�6�ե�0p�Ky����Z�KK�u�%;��2¢s|*����d���v�������+�����8^O�^W^ν��
��]l$�U�bJ�Á���@U>>�m�.<��򪪄����Xo ���Y�o�j=�s�kЃ�%a��P���c'ēfP��
��=3=��;Z��:�{���_5p�3.**
Ԧ�j��=�5���̹�9{2�2jxl�_�HO���}2���x��Z���Ne�mieUU�n�\�]>�u(.&�I�G�Ml�Z��4�4BZ-�	4z��]F̆�r����=�sm49�ri�Y��-K�̤�$��'_Qw{7�|����su����I���ߠ�'�����aq���p�1��'RKdو����ɢ��$:1����d��N���uȿ�2:BY�.���5A��v��@�g�8�H�#�ʶ��[H@�M""��,)��XW�v/�꥛d\JPO��s�_��W�s!e�f�"e��n@�[h���;|�ZXǇ���߯i2��M�����ӿ��P��1H;Ar�I~��aZ���|��ȰϼP��+<}�	���aziV}1���.����g�ͧl;H��C��VGloKy�1��h��7Mfk�M�JxO����z͎��=^���y��R�g��Cf5� >8$�ٟ��2��<3.�O��%���zdE��G�M7₇��ԔW&ڔC���2�:e�<��ؕo����X8"m{��(�u%�����Ur�A�Rd�f1*���e����A[=����b<+�/��Kt["�ŏKo.�3��}.O��,��GΠ��V/����ٙ�;+~���5�y���T��?�	>���Q�����%��,Td36i�φ��^�eIrT�'E5�-d�8,Q�c�Y��2�3�����P�9Trh}�i-��~�Y�T ����T=7��:֓��z���i -o�(7D�?���P}*>�o�t�U�<�E�mU��m����)�:?�=�����f#���g����d谣n~.�u�~��wش�3��6jGȉC9��̸������f>�����D��w�������GvKF��W2\V����DM��$�"8�A{��qm��g(D~Va��|��� s�*&0�q�c���E�Еz�2��٦١J9fᣌ> ��*~f��'0��ʘ��n}��9ߟ��傘A4��e�Y$�U�S�����z�h���dW�Pi�8�Wr�ɍ�]")\��"]�R�t��Y���ʎv��\�L�Xx]����4Џ2h��¾�^s�z6�������À�ܧ��,�
�~��z�m��/��Ѐ���ݧT�/*�XkSd�|���4	��GfwRφ>��a!TX��R�}$}𙃁z�O[ L��z���HP�;�C�����;������,�)_'O�, >����~���ߣ�~DL>�{m3��וo8�`�W"1��,\���ؘu��Ԃ��������F?eg�$g���=�&,��7P�M��?��̖��S+�-ҷ�u�qq�t/��gv���ɬ�[�a�j�1�I���C9*������P}�3X�7�����'��[k�h���B^�������T������*m����s(�[R�x:=�W�p�@����w���B,Y�`�
��+c�@3��fO����;�����aZ��΍����=�ڎ��3�* +쳁yJ�71D���&�!�̳�孔Ϝ$ߓ���{�k��(��Q�����;�-d��+j6�Bʇ�Kzd�8�%{q(�N�M�q��k8�nh)䟰		�Yز�n�{�j�����J]{���ohĢK�0w%t�_�E=�W�ѯ(��/�8��檭���Y����ڊ��.��t(��d*�<>��5Ө�a�A�� Z�[&�4�����c� �����J�%2�8��C<����ҝEHS#�j����Y ��֢�U#a56
� ^��l�~"�l�g3~��Da!�g���e��6��T�"A��[y��s�(���d�I�P��d:�a�!N�,�̀g�J���q{�!��H�9r��g��,G�0g�t�ȏ|��Ίh�p�$���6�qɅ⾖��ga��.
 -�f���p���ɍ@,��rv��:�����H����fY�h�8.��Yҏ�ͦ̑�u����L�?�~�U�C��R��R��ox�[	0�4o����8;s��B����<eZ���C����"���p��w,��ts��}�\>�ΐK�s��i㘘���f�o�4(���6�:��>Ж�J�����HX��y`�� 6�)ّ��]:�M\�'fJ[�9\�D��\����t'雷�:#���k���Rh`���V�I�d����e
��k��Y�B#�+������$��+�d��G�47�-|GA+SP��H1=�bݤ��ן�l�L�&�/�yl_ߕ�b�u^8k��� ��R�N��Tm}�l)ƶ��==���}<y�xt^���@lq����q8�B�M2����Y���tX��]{�/j��;n�c
z�7lX{�bcM��@yKڰ%��@R{�9!1kgJ2S7һ���I7:V�p�>8�S�����\�vZ!�2�WF%�g��֦�(MҹdT�t3Z�����<!%'���.��_�l���B�G϶��
���[�w��$1=7��;�׸d��2�$��"5��6xu �1���D g���S_��Lުy|c�{''��~�)8��_?h�6F�ڢI�O@������GSx%΄F:|u{+$�0e�m�a8w<�92���%2����������[,��hWg�����E�[7���}�N��z,��ѢZ[��T�ö0���M%���'[�w��v�H��s���R�b��`8��kɏ�*$�1*}ֵW�϶L&i������|-^❖��#�f��.�UuF@�� ���$����v���()��g�U#|�ߜ\��V��7'���U�Խc+6�Fʡ�(��Y�ׯ�G��	/�Q5��G٤maD:�P�R���\��d��=���,̵)�7�M\�+ʹ����1�@���#/��<�X൶��ׁہ�p��;�5�Rآ���#����Z�_X��b�w���J�Fߪ�VRۃ}yG}���[n<]5[h7ĉ�EӺR�d�1�jw%޲�b�q���S�T�+�0�yW���XZ?�KI�R/��s>e��'V���Su�/�I�_.��D}�oi��6zj��9l�<ܯ�?��lA+��椬Ba��g!�OL0�xnM$ �O����d�l��9�xVJ�[r���4��݈�.��jQǭ��y���fy�*~?��k%�tFI����EN;9�|ahaA��:��`46~*^�9m�V�gǞ%��JRR�h����M���|"�¥6p�j�I��<�O�w#�-�(�מp����%3��V��hq�xWj��|���.��@���T���ؒhE8��n��4��z%B�-��ʼ�O�0��u\�O���	 &햵�]�^N��=��h��΀P�$�MB뿠���'$�����C�-L4f�k"�*��.��]�GK|�SP���MV���g�~�X��]��W��U���8*�|��A�e���ٰn7�D�%�(ɇ#A�g��������1mP ~��_��HlT$�a��p�Q�p�ԩ����-�$��{E�î����B�y�aG����8��V��Ew��
��R:����U����R�H��Aj�d��q^���~���M�_2
��]d����si<�"nV�;ك����t�;L&�H�GU�}��4�@���te9�Z#f5�P�9/2��T�Yu[\ �̖KDr�����,��K�����֭)��0?��P�7a�xLsվ��.¼.�����v����Wv�@����W�'��A����0
��y�R�>*�u `y��vR<��A�ܥ�"{i
e��T���^Q{��,a�	1�6�
�%^���ؘC��7�a`�Ҫ�. G�B���#-q`D4&�x���N�0�g�Ȯ�B��؝���**���aب��8��9����d]�3�ڮ��j�;J♮���,h�*�U�mO�s�p)O����?�:�ud��P�<�����(�Q��(M�rmx�������KYj���n�����a���������l$���u�Ӓ.�dQ���t^]4,��'�{���P	�<΢/T��m����*��!�Y#���|E�
DWG%#yh����e�_t�wyG�J�xT�K~3�`��i 3|��5� �^�LE�7RSp�L��e�r���~S�H��\mސBe&\ʿ�qY�$��h�^��Χ�k�`��F.G������&!砚�x�]�ӻ񄹎V�j�t��W�|��sm������p~A�ջ�����
4Pt�n:��fu�j|#w8�A�x���'w+8�i��+:D�U�u84��q�_If8٥Jβ�rÄ!Y�%��?ށ/���Ewc�BC�o�:wS"c�*Ce��	h���av�#%�o�UK:�N�������������Z)?�>�Z�����B���o�j���~�1��n��3�����i��:jpC�G��f��<�[+�]k���[�O�mE�W�HϞ���q�v4����-���>{pB����l�w���X��?�#�N�{�<���U�Tl�?�\���8e��~�-y��D8��׵�O��W��
�;�Rn�`��vs*�G����R�Һ��#�c��҈���]����`Tm�d�M�(��Nn��~�HW_]C�s�j�ɦ(����O�ۄ�O��0܎��]�F�q�n������Ec;��0aN��-��F ��Y�곮�v���$M�*�w?-oի0���U�|:q��g�Ib�㷓m�>�z^��j���A's����1ۭhݶ��]���X;b�@��%�->n{!zvh��R��@��T��3$`�tgfNG
��W�wO���C:�Z�tL0��n=��Y!4ғ�m﹨jS��!��b.Y��P��kQ�%/>�V���F����8_%�5�7� ��d��*�j~ִ�j�e��*x|����(T�Ŭ�0s5T���psz��u�6��Xڙ�H?%v͌4Ū���-ߜ@v���g�nI�]*�P�%�m8v�DFJ1�Jm��?��AMY� �����H���cX:���G�Q�<�������2f�PK   �}rZ������  ��  /   images/a4634dc7-be5e-40a8-852b-d0b700abe16e.png�{�?�o�7RY��
��B��,3������=Y!dd��:B({��d�!;۱�v_�����p��y���xw�5^�9�s��TW�EDG���sKEY�9ε��	n�'��h�_���88ʦ���{D~��O}OmkO/3w+///^;g3W+^w��MI:fyY��)o��i5������d�����N��*�a�U7E�����؇�x$�Rtzܵ��l�)�c)���=�n{��E��N,�Q�r��M	ِǹ�S�=��nF|P�26��������8���{��bB"�{q=��#���~���e9��^H<Ձ���"qn{�����o%��魡\wq -։ov�P9���ߘ	Xz*�p�9��n,rcn_9�"�I��K���nɒG�m]���_P�2F+h�2L�������Tm|��u������Q�7�Gù�^���]�,sD D�S����L�Z)F�0d ��
yh�Q@Y퐛�\|�E��-�,���A��Ɍ��;�(|�/��}$�������"D]^��N���c%���?�V�7�+�V���fU|~��$k�/�o`c�ԭY�`�R�u�1���Ѵ�K~��c_���=`⻚�͌��l*+A�n���'BO�6�+m��;F���M匡s��~9�󭒼��6ꅛ�ˍ����C��lJ�	<p���� /pkK�M)�b�ד�V3���666^�a�B�(��B�KII�s%�-�mB;ݨ�C������*S�����O��*hM^��.ƹ��pb/��]DDٿ����Fk�7蒇.�$ח��0<�%H�yבJ<�	S7��pOe���G{ez���3���5n���@e�����'���V���p}���xU��ߖ���'PD��� nI6Y>��{v;�t	B\����R�Wk
y-���Z�C��NF$6k,>�B ���ة���ۈ��Ѝ��$g��8��s5��8��S�F!�פ�&��+'�@-w0`�C��9W�W^���-�8��<���2>�˒�P��%�f?�o����{j��_��U��-�ϷC�G`� �s�8�O;tBXp�x	�zb��8)�]\���RB #�jX(�1�6+��­!n�l=O���#�������%P4h����"(�׮>���EJ�W��{�.(ϋ����y��y"\6��<� )����������b����9�r�Lp�.n������4��|�D
�lO��8׸G��H����Y_��aO�~�%8�L�S��P�v�%\�cע̾��!]��oNf�E0!
8�U�e��6p&�?�	�X-x��>��c2�)C�_~����|�O}�~8��K��	O�~ɽ_�]E���Jf�*[��@�TN��7�V����˒�����$
˪=۬��g�,��K��{�22j��5�gwp�7�K��f����G���8�4�l�8Mh��4�z�]�[�&��T��C�I>9��t�ߪ(ˌ�:ѭiL�3Yp�F�n��]�VR*č�y�+��yQ�uY�k�iO;=��it��+�!��T��N�Z0�#NJ��>����<Q���^�~����y�BJ���lKc�Xʎ�,z^T�$L.S�R]�7m�ې����G���3����HOUԈ����#c��#��9�+��[M���������~=jڹ��V\vbe`��F���Y�|�KT&���;�X�W#t�s�v���bӋu��U����޺X�G�֐�؇����h;���i��q��B8��Hc�t*������zAu'��_�ޝ2X�#�c�`?�ԛ�kӗq"����W���Q0�9O��vy�d$�^��˘&  �՘&���"2#R�$s�<x�qu]9��t�d���Í���˽�إ���x{;�d�X
u�,���,?���&�q��4A��.�s�O�So(�a����*���3��2��v��|���3���]W\�]�m�F�ި�ݼq�%m�Օ�]o(j.�R�dV�{�&(ܓ OZI~#9J��������b�w_�Z
FZ
�>�a;�\��Ml�rc�?80��Na�&G5����<!k\s�@��m���Ro��ׯ�,i;�0u�yG�*	�vCl����B�@vL�i�Q��2����E����W��/F�a��"�kH�n���X�j7�]���Df�\v���>Q�r��wT��p�������XN?{b������bώ�<%�%}*(X֝����G�ӳ{�m/ɨ$�ٴdC/���	�j�������&cs������^L޳������2'�6'sI����൉2���?��ق��G���/�����n-��W^�d�8)g�]��9�,����U���FA�)��úR������ވvs՟��-����"�<�!�w��� 
��b�}��@�`�RH���w(v������p��9irH�%�`�K�H[��f�3�7ov�����z��+5�s�5�c������lS^w�W�&k�"A�K�71L���3H��գ*�Z�C&�[W�
���v�b@���n�%۩& t�-F�@��-��B��R����b^�3T�筭�Z�S! ������v�WS����(�g�6h+�oC�ɱY��;��t��0�����*a~Ǿ8��Z�"�dc@(ż�Vcb!�C��$45���cۭ �	K ْ�������"�[%<���,���Z�<n��C���q�i��7~r9e߫�+�!�d؈$�Frd���F���Y�ޒ������U� �Dا��J
�s9�l6_]��53C��b�ra0_-��wy�
i�g�|�W�RA��z~�z�;��OBIt}����b�.3Z��p��2��=_���-��W(��pwz	HR?I!2�\�j�������F����@Y(B���
���C�"ǌ�Z4��m>�i��G��汪[jß���3���)��.��������X������v�1Z�Y/�E	����D�-��z�#��]�hc�2���'m�j��Z�U�3��q�.��E��A���d+YnJ"Y-J�\-���|oT;t�D���h�(��v��n�ݞb�A�FZ�VV]yB�9��U\	�ھG���r/%$�\�wE�iε������k-�ZP������s_���ۑ5QJ��1��U��`��:�]�Ǆ����Ӽ|������ ^l[�����W��F��6�)�jqF���2�	GD���!
��4&��i�V���5���&������9Y���_�U�SM��O�m�⤈�'nz����ۮ�&�l0���3jw6�hʋ�+1 a1����vb\"�ix���r��:	ybs��UE.�ž���Q�3����jw�~�r�|	�xM�	`Gq������n6�N�S�S�d�!�"%,��QsF �z�;��	� F������6�2�հM��)<j�/YO����"���rK�^0��+���un�_]��t� w�Ŷ6(�I�F�e'Xvާ���cz�0�DU|���SЙ�9����e����D:LMM����O��q����"*C���\Y�FߐI_<�8y������Z���h�[3"�@��xe�su�}�d+���}�S��R�-����p&�ٳ����;�ϩ�?k.B���:ڤ�F!k��Z���sJOk���2� �"���L�I��,(�BgP�:<�ٿ�	3ш���<7d�ϳ�"
ykK���`�s��^j�V>�U�=A'��CDXt.��֛.�P*@"�	�J=`�ce�{(���rc(D�`.��x�
'�l*��..d��%!��X�.Le�6|9"ԛ:��i.�FAa�6�O�Ҽ��/:'�p�=�B���䜫~L缩�v��G��b�3R�N��j��g<�D,�ꬔD'�|���e6 �,=��x��9~K��l*ar4�[�R�N����
�����V�j���b�ho  ��f�#7b�%'�n��[Sb��Cwz��h����1Y�]�D��x����<4�1�ҙ��`�2[����b��5�ib ~�����o�]i�n
Yx�7ކ�ń���]h8�K/�L9ءD����hH�,Ԁҳ@��yL{p�56٧�Dgי����iy\'���<W$�.��7G�1o���a�N7 �x㇌��=���4p�Pٿ�bn�n�H�/+^��t�hH~�>]���pՓ�m�:�绽h�鸹9�w12��CO��iNL�S�R8�v=O,��6�&��V��_�>ϡ�r�a���^�)��L�*����5��j�2B+��'�9A&��A��w��(���.�X�.����$��G0��:���w�O�/ϒ�.Ҵ�� rF�U�-� Dx���ŋ`��:�a��nK~Q�Uv�ƶNE|.Չ�4���`p��h��Uv�'��Ug>0�
=ڜ�X�2�s}��վ��S�m��l��?�� �*��U���䥭m���B�d+3o�#�kQ��o��~4^,l�B�X�D�����h�&*�|3� 
	���*h��%�����J�Ak)h���?-�|P�LŸc*�aG��G���#@�#��W��*�?��RȰ����kjÌn��R�xe�n��ٕ(��`�l��}�J�e���=837\����4��p�$�	>�D��
莞�g!��D�>D�����	��Ӽ5S=pP?*x����Ȟ��;�`��V�jJ�U��45I�ܺg@��R�'Z�x�24�������"��aӦ���� H?yq�u�V(�R�{D�TsЖ���*��韈V�b94��.Җ,VO����TIX�$�m��&���:P�p��G.���>�bjÛ�� N��IOYH��F�t���k����+~o����<15��jo-l��V �FU9�.��ǭ�2���7�&�m�+�[ĂB�����r�4�R)�w�qPW����Jj�_���u����m ���{�U��ݘ�0��j1+F�/L�́�3���u��7[U�ɚ�f`cd�:S.��P�Z��c��#E��1UUUH�_��03�x�~@_y0ך�� m�I�L@�"������|��Hx?
���A�,Cgkw"�����k�*�e�ш��1�/��nS@�qA܄��mEU���i�b���%��#9��^7O�=G�49�����N()�	�}� dKT �U!�Tn�4�yzƤI�ۚ�'�HOKs6i������Bd���y+٪�2-��o��^���.Ƽ���G�FyO^c�4aT����B5y��TNo���g�<���5�5��e�.P�q'tH�z,�~�q �bPT��'�l�NY ���6B<�{y]5!�W#e6@'�z��5� �Tھ����.D9O�¨�]�Z����˩/����.��r��W�W���O�IY�uxn Mb����>2�Tࠎ���̮���@Y���D��Іv`C�;���4�x�ji� �Q:; ��O˂f%�2�3��޾��m�?�ܛ�"2ꇀ�P蛛dr�ߢ�����v]�{M�7�)�49�#_��߆db��NJ�����H,���PfB�° n$��?�J�쯋��ٙ��]���ۀz��ߪ������ܜqc`�	d �r��z �$ZFF�r�}+i�d���9zt�����Ȉ>,�6����<��8�T�t�뜧2L�]c����������YQ�7n���@�4`W,0�2v��k��Xs� ���4z�5Y@�K�lݪ�����?��  -ҥtSP1r�I<V�U�
��"�X|��{��>��A�Z�T�m�z�DF�*é�p�����N��t=ޞ��Ҹܩ���L�I��vt�'����'zx��&�=�tD�鳻��Nt�4
jݗ9::�R�(�g��ҳ��l�����������>��*��M��[�/tA�mo󓠶��l�N�$�������סƢS2 �ڴ� �+�C�����T�ձ�Thm���
 8�/�wR�]�~����5��(|���Q���p7-�d�P3y�a���6��i�Ej���Yeii��8h�j��?�YB���q<Ѥ��lˇ����Զ9�a0��Y����x�'Q����� j���� h�M��c��>�.�˺���hp`�ɾVo0ɱ"n`#'���v���L_����}]�2 I�2A���Za����nb3��E���#hݛf7���d�ns�	-b�d�!�Gt1������'��_b��[\\�-��p�5��)V�C���O樧��I�6zl�/ei��W���]���e��Ls�Ľ�k�vy	����<0�ft�@D�,�����@�� @���(*aܷН(���q;M���D5�z�Ks�v� �R_f4���&7�ȿ�^�f���8=�BB=�G ���&��Y%�n�-U����4FWSG�WD�vW`��>n�Y_����-��7�p����'���'	�lK��qKK�3�UN�g�����-m'`��GS���\�A���[��	������ #3-_��@w�g*
�N��R
`�T�Φ�������<aǡ�*��\L��̱�i�{"�7"��kqR=�3�U*��F��/>�� `�X�ҳ��y��5ϋ����ŕ$'Dw�-�d��f �_t��D�Kߏ�Ԣp���!6|��
��u���g��4�������κH��2@�M`sB�������9��hS2�-HL`���3�<?ib�qe�	:�p�/��t��GU�0��>	I�w^34�v��|#���u[�����F!����ы*��V&�hF��OB�H�d�����Z$�齈�j���ŊN�<����)H\"-��>IRY��:ފq�_�2��^�aeu
0[��=_].�rGU�𿻷�G�	��9A����;��k:3K �7IZr��רվ��޳��4�4�W�ì�N?�Ko���+�U\]^�.0�6#O�t��NWr�r4m�h�l� �-��&X�gŌ���,ݒ���10������m�~��WL�XP�ښ�1�]���1�4VI�����.��S|�ɒ�<��Ė�:�QG�-�b��������_ŬE0�Jx񲫦�Nd`��%��=��ܲ�bF�ީz/ uSN
�R�#srXDc�G%A͊R=:�';������h�v2�w�K_y�T@�T*i���3�O)~�?"��ٳY����t)��Y�������'���c�6dX������.�*���q0�A�/�� ��q+l�?S�9�L�J��KQD2g���X�^��$����9NT��x|��Ƃ�����nւ(�t�����&h��^�^N��Ο�@���H�)�G�k]À�)��pWw�"8��(T�V i�c��t	���ٗ)�cR�8EON�+.k���I�J�]��X|�U����rF!聩� ��꯶���H�pa__�̈І�O2�]���uvN���W?\`�J��c4�!�va��`�X;��Ecy��U0�%������׿Ňb��;Xɂ�_,x ����K����}u�4�$W�����i(�Y����ȫ���y*O@�U_���03��{l��n�{[kt��uuuM��5����������<Lx���^Ui�V�^�NL���7;�~+����j�����١�㪯vUxqjZK���?w���@���d:e�e2��Q���s	c�Ժ�����}t`�%�	�]���..�C��xwN�4�
��Z��Zo�Ue�+�B�>��`{���L�B��c1��*J��y_	^Z[{��������tv'ی��F<$S�gגǤa,��M����8���L@e�:�;�����֧��y�Kt�ޜ(LҤ��,���_x;�U�S?GT�~��v=�K�hqsu%�j:���QH����q2z��L��s�D�Hʔֈ5#==��E�e`����@�U Nl#�Q�{����q�m!ox�����ө���;��)�Fr���W��B�qR�c|���7�����Vnlj��@>R��,�P=��,��"��҂S�4�� %d��m�;:�1�)�*0C�����dq�B�34���D�H�؉ر�T�K�fK����/!�DG�k��XH�Q��K��xY�A���E��4���GRc���,u���p���e֕�q�$x���9*rM���a�"ϣ�a�SRQ|��� ��w%^}���ɖ���X}r?��a��1�,`����d�d	��C�''=T�T�2�"R`*�C��t�ê�
�����f&��6*�l�0=�v߻�9��������H��ݭ@�W`*���`觭}��9WZ f�0��v<J�y`n��3�~��f�疔�Df��vH�B`�Ą�"�,B�u8�*
,Ŝ��t�''S�C!2(����tC�	_��9P	���Ҋ
:Y���ʰ�p�#�y�.QG)d��(CZ��o@����7�Mq	��/v�b��pQ���y�YF�jy v�-n����A�S�4Y >{K;RI�<=��μ��a#q^����qf�0�RH��w�j!}��;!��zߩ�9�C="���s�l�|k�l6�k������[ɸ�;�$v�HVߏJo7�VV��:�F�0�
ĭ�ڰ���&;�9.2c <��w�m͘��i )~�1�c��,,��M��1��g���pc+��B��
A���59�숛$�}������,�x���̣�����פ�)3��#�=4�p�>�Ӡ��CI����7���XY��u��"ʁ(.����Km8�㭒009I����.j�X����%���{_ ��]t[�n��o���4bbE�>��i�`����d�P�;�Ա����R�6�'nB����#(K��w�د�N1��-6��͡>��Y���j��`gD��ɇ�W� $��Ո=�D�MM]( ��XWZ��:��c�vQ�z�����i2�3Z.���j{!�UNz�_��7뷒�,n`4UΕ���ΊA.�N@�\W���Ր�(.(X�t��i"K�HA˒[x������,�~������N`�N���%^��C�m�ni�P����3�>I�U~~���\[��}��ԯu�[ϸ����*���j��!����� _�r�[��è䢇�<%�e�Y%�����K��*�)*���ׅ�����R1#B����j�_<�)�6���=	))B����%^�,�M�`�� DQ
��>���g"���v��n�@r���vs/`��+��!�3��`����f"�S�U����;�|@E������N�况���Lc?==u�:s� ��f�L�Sy�)�\mޘx��[8<f�#�>P���Q�BM�<�U��>��˝&�*�P�\����e�J�h�>�K��n���O�-�(�����{'���ۂY�bIO(xL��_�I�(Oi%؄��`���}�����0q��B�kȃ��՚������Q)2�5�M<4�,�yo��͸S�f?�:8,Bt�(s�]D	�]w"GnQQ��L�	0DI�z�������L2�:�	~Nm2���u[��]#�t��<��8�;_-�Ckk+*�.�H0�33C��='''���^y{Ӻ4���#t{Ł=P�e��=`T1Q�!�v���-3��P�^
IƳf�5ilV��0�'i+T�|@�W�x�����;2���|��v_�&���ܪ��b\��@�<y�$��>5w��#���h�'&��%�L�H�^鮞�E�f�S�����d���/%�5�.*xK��V3�K�͌���=��M�p�m��p����3�]O�bE�RN�%, �n��	Uj\,�[��,Uc�F�~}|�=�L�mqOE�А��A����Ζ���x桿�P/!�����LWD�@b9��^�Ewĥ3�Y�bN�P��j4k%��`����;ڄ(a�>��|'䊝�%��Ũ�q�_�P\����WF�fhYb�#�x4o����q�@w=����H���V�b|[W`�	l����V�@X��eId��͟�p��G��1�l�h	-�H�d^㵢��|;o 0�*h�AN�]��f�^��̋Я��8 n��3���nP�t��pZ�
�ѝ���-))��f��*-L��J�~	윴�|�<��.�?O�p�>�������W��"��æ眔�Le2)��w�'�y����!W]À
8f�:� �|�-c4���
i_5|�/b6ز���؃	o+%�ˆ�ً�F`�0��j���0�O<<*�4�@�I��@�K�i�'5 �| ����kpxx/���yѬͿ�ϋ>̘i���ׯr�XP���*��~�Z�����^����l�O��^{��{_l�=�e��I��B����c����d�%��w�O@��q��ð����K�q�b,A�-�,�sF�"8�J l'��A�ob��%QC�����;�� ��b�����5��/ָ�$=�t���P&���ŰP9p'd�'ic<s��P}�b��{G�]�ޗ)�U�.7�%;�g����}�����˥7�8dHn�j�'Ѱx��>��g���I6�@�D}�E/��qB�>-�`�� y���?u��|X��Jx,� A�ۊ"��5[�a�������*i��{[��Kz���h�r��P��!EP��=�.K�����G�[j�Ϲ���YK�o������������Ma1�09��}�4�GB��<g[�H+i �9U_�5M��l����9
qh�F�8�;��&K}�/��p�5;l.��w��8����P�t�� O4�dBg���p)B{|hUH�#	O��̹t��uٱ/��;6Utd�]�	�l��C�={�$s���J��>��ٕ�\i%c!5��9Vu�1, �a\;��F�{�C�����ʵgDй^���GF�{QoM�r����1�����E���z[�h���y�~�E�۷=S�:���HzG(�c��	5�{��
�������wT 2:bް��+ܲߜ�Mu3�F�����h�=��2��d)�&c�(0�]�s��3L�b]�&��r��]%�q[����-���6��?:��i�5]PV=k�=g݉��
  ��pN�d+,w��v��T;g�QB��@�����񦜽Fg7�����P�"w���}Ĺ@=;3H��	.D�Z��,��$}w��.Y�P�ZH��y���/��;�n��-��N�"����D��܁���{}Fg]�p���Ғ���||"V���W�2o��@=�����ZD�V�~�K�F�*�����8� ��u�����U�����@i%7'v.��A<��V�튪o���n�� gZ�2�4X��H��;L@�M+����F{��T��xK�k�F:7��e�y��y=+H��ZP���;*�����rY�J��˞�@�����z=��hrZ*�ب�X��"�OLNVVVj� O���X㕏�R�kQ������:A;�=ޙǕ��a�c�Y'I��
��N���@F�y�y������c� �2���Dn��z6}n��7�,:�b��a]G>��:�gUZ��#�i4�]>Y	��1P��_�6�'F<oo�@j���O9�3�(~�H��k�C��?C���pӥ�]=CT഑��۶YJ�hc��ۻ����M7�$xK39�-�-�UWZ���OK�69⊍�٥y/&�}u_�Y�I�~����^P+�;��)w�	~��7.���d*���~���X1�IU���c|@Id�-(�@�[[�q�w���i����2���眬0�q�۾��1�[��К巧��R��cR����������ang�i���]�Ǧ4�������QX] QU<rVߟ-�� �`��'� �N'�����&�w����כ��|�Da[>'>�l����_�ԛ�)���<Ժ���z��׋����Ӏ0.�$��Hß�05�}˞�z ��7t�"����:�\�g�59CA����6�����������`X�E�Ӯ�� �"���pC嗁���=I\3�y�%�E989i�~Y�=�z3Ers{5Vi������ycJ�]� 86�{g.�G�1e�rE%C!�F���3���T�F/�Rj�䎻����^�E���Q�g���*'oq9������́�8r���s��ZV��2��eT@�&z��g�r�K��t뽶��pg���;�PѼ�5_�N����E��y���㮊�T�e���ǽg�c���<���~YFڵ&��Z�-W�~���ի�Ai��9�{B��{�ݼ|�(NS�e���g�]m�2v�n��5=j�D+l�8`�����}�_7_ʒf��E(]���3}�}���b��)i��Т���^�kz�������y�L^a��)h|�2�2�*�r|�:���DM��������cJ���ƾ��&���چ߁�r�v�Y�9�s�E��q~7�d�?����0{�v=ٽ�	��r[k��_oF3(wG��+eo��Y (���)�k���E+��'8�����L���}}}.'�L~&'P�5(�w3G�"�D@H�ޥ�TI���&�"BȌ(/���]z�z���4_�|j���{���r�u�M}�u�1����{ȝ�C[��ސ�F�;ƃ[Jb�A{���#p��k���"�z��Q�����N�r^��oa�og���vc(X0�%�^�2ꇲB&'Sk�����Ja�?��y<�QV�\�'�"�hb�_���g������;#���/KS]@p�\	�u��G��vK�3��h�߀�П��J~u2�Y-��E"�)`����]Q�@54\�lxxU(�Mk������:�n�"O����a���ߨ����|,���;\�0H9Y�5U�T;��Hl��.a�Dc�?T�EJ>�͹���;�|�*TIN+'''�3-��yJv�����FUi!@K�<�uJ9��%�r6��r!jĞX��s�ZaP�\D7U��w�����o��o�g�֟�}'����D �����-��^Ҍ����D�ro���K����y����Eʘa!'쉈�?ida(�]/��)$2��gL���*Ğ��.�d�%���?�se����[����a$��.�䖘��6�5շ��r:��]S[�J2>�l�L�Fs�?Sz���ʈ�x,$O�9�n��a�v�T__�u(Ɔxێ��uSJJ�����)�@귩�T�����YSjHCxZ���/M6��W&�t�����? -F�^��k$�.÷�$ǿ;�D��_g�O�f5H�*s�H�&=��^�}Iۡ'}�ٟ{�$8�8�_���j��K�֡RT[9y�uYrI�K���p6�Pj��k��/�V�K]Ц����}0A�o"JGw�
_�>��_�D�C�Ϝ��#�̒�W�S��^uϿx�B��r�~���=�m�5]��ט-Y�0m��IE��OcӿV�\I!:=y�E�l�*Ŭ���^��	�}�E^�u��U>�U��]�������՝��Xu+<�ė��\�]l���1�|�	.�� b����>��H<Aɝ��@#s�tt���j5?�ֱ�=:)� ��e�m;��aS�"u�oyS��<zhA�m�����X@�k��6���E�?Y�as=w��[2ֵƗ�K+ R1w1C�j�?�kr:f�6I���z��iȐ�z�D�PO���e�ڴ���:^_??���.�;j�k�+@�{=*:����^���(��u0U�{9a�́�������=����.-�li�]Z�&O��"ޮ�mجqgP�ޛ��Q�+&h�NxxWn#а�$��l��3���e�_�}�����ã�ɦ�w�x��}��p[��v��� *��� �xڵI_������'����Yc� )+��P�ʓ2*ۂ	�S܄ݸqc��Y�"�����t&G�J�S��DDf*��KA��\�lQA��=��$���2����i)&7B�+����f��tع�"O@���0�'�W飺|;��(@�����ޤ�il*Y^gEȺ:P\f�O����$O#�kG�bs%�ԩ�����hI����Vr���!�<%F�{ �AĆy��jXZ�<�ƣݯ��p}���2j�8��y��M�X}��U�:L?ɼ_ö�33Ȉ��W�]�L%O�B=�J����\=.��_JbF����3�A�?�f��1�(��+��C�;�_�<f��W��:tg���5�=P��y�]KWׁ�KAB��ە݄n6��P+�{1�<܂���.8��삈�T�
�ɚ2a��?=c�zdID�+�(�M��|h�x�Xp��C;A4f��Q��V���丮�Cԭq����X�����W��%�B���߽%��p��~+�U���a�����W��kQ�D��&/�%PD��;��?�����67��9�0�T�������*�@������mW5��vET�&���ͮa��8���$�ŭ�(���Z�#�D�4�&xOH%("�79�.��+v�wS�:�ڶL�Ԕ)��&E���r��5Q$��������`lW��@�����%��t{��VN4m��Ѯ'��R1Γ���;����w?�>��I}��Щ;ò���*� �<�� ��������˝��]&������H�ѝ��R�5�������N/���ߟb4f���M�H=�i2�o��Z����g��*m*)_R*j��C�?�i< ��J����0�FY��/�qJ�ﯼԆ{z���
�g�ɖ�ll���	�k:���
V��"/`���d�1�d��9�_�͌���V�a��%U�"ه������Ζ ��3SSI�,�����O�O�/;����������2�	�t'��~g���+Qk��	=򏏂U�����L�3ԥ
������|���3�y7ާ�A�}�`��G���u�o�ñ"~H��#�)�X]���y�N�ڰ?drM�� t0on}��a]iu�8/%���,�]��I���/<v�g�27��&�_�M���9ܼT�x��������NMW�ߺ����_���0�?��ի���#jM[y�8��Hޜ���|��Y�/�Wl�{�]Ҭ��YG�?�2��dj�8|�������c'o�(q�(����#ƖQ7DȠ��,��@݇�c�L��H���
`�<	��w���&nG�˱\�j����/�r�| �7T���7ǘ:r�c��_�ӓ���v	���Kٟل�,I�WJp,���a#�h�"�q��2:�4<^��i�]�Xֵ�K���VyE��Tr�1��H�o��דM5��ϧT1�������g���uW���`i�qч���<�%�F&݌[���ۧ�h�'	H�@�_ٌ!ԚBX˘��Z�`|�B�e7��VH��?�0�R�-�Z�g��|���=�������@G������`|O�r���B���/��Ŝ0���н����X�X�_�����@�<��e���C�Ԣ���/xI������!L��|�+V�ieD_����IHo���3tv|�d�9C���Z-y{B�O0i�y��+w��+MiVТd_ѡ},�����D�8��Q��&�ӓ��K��s�6�v[�q��Nq��E�����A����vb��2}O���*w*����weǼ�����67�81��f�.c����Wf5������b�-n�u}7;8�<�rG�E��u,#S��ٯ4:��@���a��Q�8�=��5����S���,:jl*r��|>���rR���T���"�@���G"y�ÍD�����N�?����+�Ա"Z��!ޑ�YK���"�F�Nu히�Tӯq%LKvȾ��iQ
X���:*�7+�H���Ew޴F~/�ы�!?�f�r���{������7���3�Qq}]]�7空��tZ���{���j�&fx����u��/��b��R��!�BBB�gU*L������J;t uImj�F� ��J3�׍�$�z�Um���ӻG�T|�t�EgdD�uڥ��V#F�� �QT�H�e8�\�<H$����	�-T8'�������*	YX��9�1��V��c�*I}0���"��R1((p(����������Z�k��;����p=K�6yN�;h�Ƶu��]�=���J[����k	 �����wB�^t����u����U,RȄ1��z&rP9g�9�55���\���!#�kMOX�X���a������g"?�ll|��%5J�T����ˌ�r4]S-KܣW�5v*�A��l�3Tŧ��v����{�O;&liж�^2����0���r��\cP���!HH��"���\]���>4�"G?��s�Fn��`�m���"{�o]����A������):�v�E5G���/��\�ȇ���������|�)j3�D/k��I�|��p�n�[s�
�y�c>�I���֗�)^��g8P� *�p�oܾ��Q�i�� �� �Ϟ,��EYj�	��=�O��y��B/��ʻ�}׾���m�܁U81d��ɨ��[�z�@�0?Dc3�4���0�㓽�Rʢ�a��7<�'��+A�v�n{��b����}��[K�2>�"ޥ�ѭ��j��%_ڝ&��?��;�-��qi[���V�JmiyOس���6�u:>���������-���t�he]�U7���Y����N&7g�S���l��:��崏�Zś�u?�U=;��@˔����
�2^��I�K�j����ae<�sX�l���AH�M��#��QjE��$��� �����~�H���n��'��#R�o��^Rj�ge+=��I�����{�z��޴Hk���$ü��6WS����)?o*���VZ@�ʍ��x��m/-6o���(Ϥ[0�Hˏ�+X����n�]�I�i�g5ߓ�>�2��F��f����?ԝ8:hH�&��1�9l�W�X_\�S�u�?�S��jl�^�і��\W1���E��n?�^Q(C��u����L���d����d[F�2��\�w����e�qM�t�v��8m�+�g�/�8Ԫ!Z둎�G+�DD8��5��y|0�νD=����K~��O��#�=̠�^k�)������><���i�n6�O}c��<ű�(˾�d&�*�1�wg�/�<�F=�S?#��Z�|ez�̆@t����ח)�Z���KCr�� ��3��E�'���������O.֗���JH��uJ��^�L�O�X	�(H2z�v�{�e��Q{29(���gA����Ƀd+�>#..�1�X���kL�����P��4H� ��0��aQn���ҍ"�4"H� %� J��tw)��tw� !-�H� �)C���<���r��9��{�Z�س�m�"���_:43n�j>�Ѽ�	I���3�J��Ʈ�;!CY�o��<���e��U� �(<C�� ?�
A�,:V���<��b6�Z��St����gm	WO����}�t9�4,����X~E��GZ�1�p�4��墙?����O�Y�}�_���3ͣ�TE����ÒED⌱�'�B`ƹ|iXA��[3��=��\� ��I�?���T�\�4%�B�ҘG�A��D��Ʌ�u�\��"�	��)#q�_Z����:]vt٬�������˒�}o�I��qۄ)��4�>�,��F���Ԏ[J6X���@d�s�+�ծ%��0$�	Шkn�`)�0ţ{������t/~��H�y5�L��2)%�|�P�J�e���A��uϓ��Id�����a�<6I�?��/H8+�=�ۍ0»�N$Q^̤ׇ@��<ߴ�4��o��w����Z=<��e$�OG&�(���jSt�;V��C��_��p.K:t����Ȟ�_A����*)f�\��*�S_�Ϗ1z�ΦԔ$%���վ�fO��Orɿ �Bo�V���l�V0���&p�MO��o#�y~V^xh8�Vu�]����V���W�+G�ۨ�7�l����+����Wl�X�E>��5�5����ˑV�T��/�g-���ի���.r�T,f�Z��lW��_pK� 	򳧔ύ鲩f��r�~�)�IѼk%k���ȁE:X�� �d9��=��N
V]�3�~{1���9���N ���V4�7p���丗�n�Ub��9�ٚ��Qr���_���sΘ��i(�d�r��?�8�z7ܘ+q����/߂B>�z����%�d_�DK���Ro��؞��ѝ-F�i?��{��3���V����I����Y9no��byp�A���s$,�y�tȘ�*��8�����M>^��A!�u���g��)��d�x'�Lg��H_�z�^�h�ߔ���#��f�r̒�)����(7��ŝ�Ni��r'��j��۾��Q��gݡ�1l�醗�w�:���ѷ3(���=��%���[���H����Q~�i���>'d���ab[2&!dw�[D�0os�$'�K���`ц�_�>ÜN�e]�_v.(0D��?^OT�����|u�'�@o�6y5��J+y�>�iw�f���G��E�����5�0�\�
7S�@_��O�vZ��&\7�b�ݜ����L��b�[�i�3�u�Y-xV��ߊUua�@�¥�0��w/��1�	�\f�ݭ����݆W	8t�/�}+�o�%1}rq�L6#((P�:��F��I�$-��8���q�O�Ӷ�H��%�m���#J�2L��%TUc�dfm��:��Yx|_���2�;h�2F�C��bcNOO��*�
0�8ѳ8Y;4[&�!��of�!I�ML!�e?�n���#��.��G~���M���`���_sM�s�'.��d�x�� D��n��w�N+ t��.��hY�)��M��L6y�=�&��օ?�K�+'
 ���f���`��JTʿ��X���=�!���IG<�I���Q�߀���MֹHr9<���-\竇�l�(���0����أŪ�u��7�����#�ZCK�JT�'&cC�{����oR�ѵUk���P���;)�HQ��:ʂD..�w&�=+�a]Xt篤����d�92�F
8H�m�����_���c��Q����	��g��P=�!Ò��%�G�V�hh��}?������6��/&n�jNI[���"ə�Tp����c�Wb��߭5gBU222`]#�s�Z�]�Ex�<�]�7���PJ
��.��)1�)��ۻ;����"�~��B��\T�S�BR��p��ֺ�'ى���
0O���#2?v������]ݝ�۠�[�P��� �b�xV}��Y���㔚�{��k�����h2AZ��tX'`�FVE�AWz�F�GjM�C �<� �X�c�Wzǽ���8��6|�%��M�Y�7�4�JY��e����j(��a�b���F'E���C�Z���?��E@)��bW��ɽ*C��d��w5���I��=Sc��ii����!XT���4�`�����r��'��*��=O��7�E/�^?a�kN��~�5���h4~��̈+�-U��:��rw�4��`N���a�-���qs��YpJ�˷�hTm��~L�׫J��)��C�54�>d�ښQ�#���p�-��qDh�v`��4�|��Zx�_�o�<(ǆ�8
3l���xS�O��)i����딗�(W�O�Z*ب��#�d����Sb�������859�T�KyX>�Q�hX���͖2��cd��=�����5��6��Sl�'A��XE<I�	jK�����|@����I�DМ��t��IJ�2�Ԉ�c��R��)q��p�������ok����E,���̱�M�?.}��k��^�bRܦ�5���>��
�^,***|��a��A~�Xt�d�R#^?�]f�$dD����O�=�pS�.�f���J�WܑI)��f�~��?�v]�����owJ�c�g�_�f���-J�D5�t��>M��F��?�NN�?Pt�B�o�R��c!|�pNBB�RK�Q�߈K�I��,3�a�4���Ԯ:JKU�?3�."�fh��twg�0MG����X
m&m4r�f���v���Ѷ��^k�|-�s.�S�y5	�7R�%����[*|��@D~|�jkޚ2 ��gR1�@���^�@H2�C+C�]�� ]TQ?�[�m�8�[2�{�`���V:�]�B�|#f����޷�F���5�5�k[��LB�J�\1aWy�<�?��-H����x��MS\D�2?Ճb��?����8����</�}ʻ�jʂ3z��G]�O���.����M*��i?����pX�hP_���_YQ����:LAa�-n"��Zu"N��{���H�
�gtm �z��gg/���V��yj2Y�[�;��~�GGG�h�\%�G�.;���e�����1�\�Cw���K��MT�܊x�x��$�����+J������.�I�h�����?Oڋ���Nn�'XX.��[>��n =ƽ�o,y...��~��6t:�;<���2�Č�����	��f�ԭr�"61<q�O�X~u<�����@Y@Z+L!�{��guNBr�fW�q��꠻l�ѳ0��8��U~El�j�v����3�������W���?�H��E�p-ޭ��N� T�-P�8f�}u#]k�f1��b��9~���ݣޙ��V ���e��]6r������Ֆ��tD��+��)%�i��r*p)))j��������u䫟�|��lG��_AJ���1�J�fߔ{Z�~�R��o�f��X٭�4���F�f��u�JR�j�%��l�o:\��x�4�F<�9﫶��� ��K�s-aF;�^��S��d��օI���T��U��I��'�O\�t��)���:����'O�P.���ٯC#e�B��?���D���YJ?����*�ݾ�$>�vD��2�)��覷�M:}ȩ�o�v7W��˟>}�]7����S��o�^����i��w��U����ha�F[�@��5c�FoG�X쓽��F;��<t�ql�Y|Y���� �f�t�7�͒�}0�~ej�}��>)k���ɟ����	$�����_���DːF�o06�7�M���J�.�`��V��[[�Yt(�#�oҬ|iF&i�1�P����S7լͶtP[\ľ+�h7�����;��t~���\���6}͎_:[*[qW��^�����$����� ��i�h���;C)oo�!]j#eڄ,=�z��,�sU�hb��~���,l�Nrp��`|���*&����uKtf�$<:���U����ـgҢ�9G���8�xy��oX�s���(Ή���6V8��S�M��W�~�5]�$�b���� ��N�a�~^;��Nb�?~�#�%����#FS/���m�,�N��$t�0�`��8PFo7m���d%v��ڎ/���7GC_�E��x��ת�I���S8��Fx�.���9�E����u+o�`YENJ	����	���l�+pl:���t��ӵ���
n�ֿ�M6�zo����!*,��������+uu
��.+�fk���!</���G�W�����Q�ј?1U��,�!4��m8�<��W7�s(t�o�Q��qs�E�
����ˮ��k�K`w�b ���j�UA�9�f��|���Ã|����M������ed��MQw[�n�Ҡ㍰Ԯl=��Бy�����9VMYX|���^
�$�d�����k2H�+M�������nC�i���1�P"�/b	k�#�~}�|+  W����M ?Ǻ�SC�̒�m�����RR"�?��0��8���\�æR#�"H���J��J�۶��3���B)�s��>�d�jL�3q5xx�lP�a@�4fz����h{�*c�e�*NM�;�� �.S�>��#a��-0�Y�lf�*����*#3���xޛ%�
[�Q�\���@{���Qd=�X	����Vj�����E���vs~��������m�Q�O"{D���_Q�0�SK�(���
ķ�����uv��H,���d����UY��B./���kf�bC�'f���aK
����P�V��p�N�͊A�!��x	3AN5����2-��¶�B�:-v�ܫ'���� E�[n�*z{�C�$�a���W�`��N;S��񼰤�E����zؒI��A�^8ml@��e�f���ܓ�����À�gg-**z����2z@�SN��kEnd/MD������@z��u��G1���nls!����\Q�>|5��}\j���
�mR�Y���2���D��%M�>K��g�c¼N9�H�W�C�_t���Րhk>&L(Jbi��(zs�\�BJ<RU�����w�n�V�S	��ɷoC�m���a���R��ׯ_#�J�#O�/[9��'Ŷ6�]C:G�f�t��M�_^�w���j48Y�r_⢣���scج��%��'�=~ƀ��&kqo��9��#��.ܾ �X<�P<�:QlLS���z�P���"����SS��4�7�4�|s��4� ώ�qo..���9Wq��ںY�7�]z��C�/��4�ٔ������S*z�|Y����g�p�b�
lO����o`gggp�����DLN���f\��<�D^�=�0#u�g�J
J���zG��/x$gj�L���ϑ�V�}s�H�O0�]�_�lLAm�й��>�\�z_�f�����6K2��)�U]e��b[aaa�p�~O�*��c�;ޮ��#U1��X�_Do�VQE������������%��X���e�1��������Zy����{dTT�"f�^K6:�4u�x<��>4���{���N]}�HEw�Qz]�$���{���""!�<� ��`�,�}I,�I�~T�5xP�"$�H��L�U�j\0�gv}���-Ϻcm7��|�~��ao�	4Q�@�}g]���p)m$/��D��bE�{} y�S�t��Ī,֢K&C����R0���)t"!Cy��c�w뚍�\��#t���G`#kf��;փ�b��H���"o�]��[��pY>�Z����*gC͖v����2--~�O�ڶƋɤV�BB������c���`$�.#'J�@�����1�pcC�S��	��3��p������@'@R��m��O������x�?'��\]��J�ĢBLQk���暧�*��G��\]���,ٵ9�6/�V��]�*��	{Ӿ��Yk_,+�X* ��ON���>_0	��7RS;�< �B/q���YV���$b�wH�\<����j���� v.\���kx�V-��i�������̗�0�:W���N������4�^����� �� ���l���2tߊZ�**�������>�ɚH�<��S<�ac�n=�44�5�V�U�A�Z~�V�4r��Ql�� ��G���_���%!�]{�����[�̆����6/4�gB.��/X�O��[�v����0�|bK�f��?O��6�i�\�	���Eb��Y `��>T����PX;]������� �l`h���w F�z�2��˃�Z��
������װ&�僳���9�gZ�lx��Ci$T�-���</m�M��>{D6y�D��n��y֛�6Ǘ�����[�"��G�N��*%��\r����k9�:�;�PUQYxhe�s��������^Bb�>VV����o�<) L�9b�y{/�$ ��)�j�/�#��_��	"��!��p�3�&j 9\N���5�G�;����O�8wxBL]�6�]�s��96��Zfr��5:K�<m(���|�#z�H��7PUW_��.�8��)^���؀h!�M��$Vc���)DhP�r7���۩Z���	q?$0����H�^!���+��)H	�ľ��*�N~�Q��y���|�ڽ?��g�(7�M�O�BD�ܩ����:Ag7��>���R}��Ģ�(R����[R����Oy�Q��	�V=B��B����B�^� �7�w����MC����X�f��*2��jT�F�_"�8B��������:��*�sD��c�l�^��|�1�Đ_�$��	����H,�2�0�ʏ�_K8�ko.��U�V���N�i҄��l:L)�bҡL9gE̹�)?
��ϽfI�x=q��W���+�?��r˟,��YQ}��ݣ^=�Y�_�zh�1�M<�����g�o��(�s{�qދ�󍝈��-S�
5���Cm�? �h�,���px�X�r�EB�62%8 L��Z켫n'�����D�Cj#4���k�YK�I�������Di��֔�,����u��!2��9��|�� .��eU��%wPS����6�����Z� �Gn�O`~{�(B��j�ԕ�|��eQ�0T�󌙱��j��H^��[ĵ��ׁd^���T���5%���h.��ȭ��i���S���]��ZGW�	���i�'9r�A=b���/4_���~��䱒<�F8�l6��k�0�K<iN�0����қ������s1�U�[mƉ���A%�ϩq�Ǆ-Q�o��X�\5�JJ:�yg���t��7�9�">I��xp�V�D��m�jj�o���/�eD��U�o�	�ec��]����1#�൵�ꆕ�������P�A܄'q$�?�c��X��::8t\^\HYL�ى"�D���r�CY���9��xNO&t����Ӟb2�����%[���-`�^�]��tٝ�Es¦��֔.�z��o�]�	��z�A�,�d�Bv�~����Χ���������� ә����E��c����=�n<�:d������%V�s������pZ�p��uT.������W����^>����c��}X�d��j���/_`�㻃��u��.n�Nx��܁?��7��o:k��L<_��紼 �'z]YbŽ��Ӟ@�z�F
��g�-w@����w(X�Ű�$9_�!�cj|w2|"mN.�ϭ�b���L��}!����Hb����76�`)|�ь
m��C�e��>���!T�h�A�x(U��DxV��L��%��c�i}�L��}�`9��ȑ%�2����r����6�����j?,D�8�|��,l��켲2떊f�`b�	��9n�N@�f�jκ��dpB������/�&CYee{4���&�<��w��2�~�����_�5[�g{��s�/�0���T�M��o�b"�Ӽ|�UW�w�?I���8��?���	k�Ph}�Ȉb�R!�.-�J�fe�^�6�fO��gDs��o}�P�sT�۬�ݵ�Sy�L,�S�$h�;'�e��=��'�gckK\Aa��[������w�
C�(*b��� #�Ǥ�mb�z�	��b�l`|��|KI��yT��9�u�{������;S�e���r��������aR4�q��ך�v�,g�mc��.O�h��bΉ+�K	��z���-0|�O�����[�����[N#����"�����?�p�%'���%��YΚ����<�'ssE]�!�\�H9�T;Nxe%I=|�9�=$:�cZ)�ѧ$��-��F쬴���spr
��++)�`#?�b��}��^o=�{��7ׯU����v��L��}Ӂ*;;{L�C��	yhfV*�����W��<��4��x�J_KJ��×c�u��P�׀4Wr�����$TL�Ꮚ����fmb����������ry���H&�5���,		+*jjY���Q��/�%_&��S�|�k���y�f��*��+R}�4�L�uxjjK���t8'?��c�`>v����k��X��eks��
6���י���>ꋄ#|N�(��պ��@E*��������w��84R���6>>�?��
�F�$��P�3l�$���_>MȈF�w%~��~}0H�R��A;��n{K�r�V��Sb乊CJ"�Ŏe[-����u�:��+c~K���8�۫�4�{@��gO��V�%�7!2H
'fg�K�Z@�5�%L���ș���vS�@���/؀��s?��}�D��܁l!y�&/z����>fە�H��B]�q�8|�PEb�}�3q������3��X	H^��1ޕ��	Z(B�p�*�x��IJ��F}8�ʺG@��h�.���P�w��Ԋ�p�鎠MpӰ�͔�V��ѳ0y�+fz�斗��K�J ��������s���*R-f'!��2l�|�����xC��S(��ӮN��o���#��ȃӅ��[ ���6�Q9���*�怂3��� '��w�F�ss��1���ԙTj����MDc����54n��dT��P�T�O�&��������g/.���P$Rl@%=�!�1T:�P�Ȅ��Ssй�^�]QF����1�" 
@>*KH���I���l�Y6����9lW��E:���U��{���� ,S��gؽ'�W)ј��c�ұ=���NS4E����6�mB�+00QI<�y�-�d�_�r~���8'����φ��{`���iN���������[��J�U�[�׊�+]TT����EZJ�����Jo�3l�}Pb~A�Iº,�4P<���w���믰�_��.����iȬ��)�qF�	L���DCC�����
}>v�>倂�C[�M{+h
ظ�ۉ��p�ՓTغ���-�33)�Ap��Ƭ,���44����HɈ\$���	]1G��գ�	�j���=�|��At�ka�1,M��M������5(h#u���)�Xe�
lf���V��ӌ�g0$��Sv�2N���G�::9e54�O!E�E��	
�c�
3��wc7�a�A�cIn#:�6f"?ƭ�Bz�$�z���rc�]Ww$n��lS���f��QQ;O��GI@}�O��?ڔ^nl��A�d��]��QJLW[��A���ڬ�y�LJE��$^��g�8!��2,tTנ�}� ��[�
t�?օ5�HERe��9؋�2/t?����0�,ə�.�^��dX~�gY}�@�v�K�7d�e]]R%���2�p�Rѩ�#�|Sɍqv�Bg�X)�O~i�g& 0��-�h��X���v��OЅz3���*�Eq6�zn��!@�/LW�X�Jf���W�-��+���T��<[��'��joS
�(|�0�Wr�՞�N�@Vz`O5���rT��{���F���]�8��~�Wy��%���v��ʅgO�;	z�	Gda�:-0���Q��V�c�~}�z��?�;�0 ���݉m�����Ԉ;��d�� ���K�:��.��2�� 2^��ڀ����F�_�#R��Q�Q�7Kˍy�(@��{4���y��+?�k%ە��,�A lBכ��KDqaa+�؍3W
�݃�y����� YU{B��)'�Y��g�t�7h& %�j����g�a*��s?ݏFgi(��� ��r���yr+��QcE���|�4��RG0�k-m����Qn��`�@��MV_�Do�C���j��a:8p[#,����h�����B�n7��mWzg#�����:=����lW��}���i�>^\\l��?�Ϣ{�������e��+[:�s�=��&7�؛�ل���f�i:�2�	y� 02��8���_~��2����a�x d�k���M�H3� e�ܲ�y=3Z4ň�T�>BA���d���l��LMMEe�b��{�3���� H��)��(+էDmL��q'�������?iaK�*��w��Bdw��W�J��ű`=��RW������$����}�	0��N�3\ �\��x�(�t��J�p�L����S�C������ �
�k�eׄ�Y3f55�Uj�X�+#�9p�.V+mki�������ָG#��l9��B�^�͍5�z������
-��a�z~Y�O�9	 �� !bA����������:{��kr36�x��]Ⱥ���^|�Ղ,&�p�e�LK�a��lYL.��X~�\��A'6�Q��m�b�`A"yBq=�F�����$�J�ь�Iy����UUU�_L�콶��=aB=�g>'fcg'��D�W
�����j$A���X~�C�kF����>������ݷ��M�u���ȧ �P@�[T�&�w�  ���+@��]_b�G���kƹ;�7�
��T�$�j��g_����1zzz��*�n�yz�u���,0�!�:_�$�2�v�ܥ� ���\:�=��`
J1f���x���qƞ�r��C	�s�q���ۮ��D�o�����S�,��Z��caaa>�+>)i�#�~�,-�!��-�|P��sR���r�ѽr�nc����̻`��W�|_c�O:$q �v�&EyxJ�&C|}}���Ĵpj�xfp�3o���|LFX���fڐ���G�O��|}�g�=�=D8`݈Qo�ۿ�E�ӡG�C�*���և�==�}�-+).F^f4��߿�/�������0��~�x8��`��H������:4k�=�l*&B���i���O~c��>l�>�vN��7����l�����?|?��,�ZB�`�Oـ�q�:%�0 J�;����\�䱽,��������S��q���u����.[�S��Vc�5y)���D~ �Y�Y���~�ŋ�cE�q�{db"0-�ö5Q� ���7uu��p�� ���r��Ͱ�ÉA�M ��LT��3;a���%HP�/t/��7A<<<�^7dy|��
h�+mm��I���Z��-������[�'�&��k�M��G�gru2���
:�~upt܄5�omo�b����s�6P3Ӄ4g�:�%4�J�o����-i�ǵ���o�S��Y�ߔ�jj��&0QQ���7�TO�y�<!���z���h�H�ժ����hu��@��m��y&��EEȭOrv-��
N�d��,gFIEe��eUԽL�������R����v	]�0f�]P��W^δO8� 'o�A�ܩ(c����*�	�j�U������ٯ�\G�r��%����փ'�q����;$��FFm�ß6� ��F�a�F�N 7��:�wk��rd�P�B&(Ct��_
o����+���q�l��v�ԂN���"vkk+F}��0��(���������j˜13#�����m���3FZ�^`:�M�Y#L���A9%pO�J'����i¡sssQ3/_It>!���f�i�4�Q�k� Ѝ0@zIF�c!�D������ P���/(-UM+h��3#)���Qm	�A#�3�ܘ_�aT�CR����N�gXJ����Ȓ�LT�+ȁ����(C�<�����O)_����AY����_lG~���+q��!6)���s���P���<~Hk�K'����j�颦���|��yf 돸�B�X�����I�~�V3C	L�J}�o��c��]`
�io�u8��� �ǈk;Uk�h(X���=��J���@/��m}�F�	7�Y�e�FM3o��"7l6`UG���"�D��2 1 �`�x��?�����CF7��vrzڽW�
��d�Ё�.�5��ӕ��)�I��k�!��^jP�"K�8Kl[0	�BA�i��>�7��`9<1���Wp�i���;v�g�p
�*�hYB�[ ����b��,��K����� .b�uD�(�fza���hC	F�f�B�yU)�uW+�����ܣ��/��'ag�}�斆t����I|oh�ͻ�	��n�"Ѫ.7�$�{@��F��q���y��f��Ó�����j2�~��*��)���&4xL����T����
�����*�j�cj���]���-�'ʢ)�`�С�@3K��;N�~�Y��A�/�O�B�d%�����񊊋���C�0�ߕ;�R$ĐD��%�m���+��vQ\��0��_L�鹇��?���E��2�CA'x0P}�-����X!I��*]�u��;�"�-#%��jp�l!*Y.elLջ"��B	0���)x~��#"�V�e�p��6{Wa����=�� ����	�Śe�?Dz�W�V�o�@�A74�-6�t�;M�`@�O��%�D���s2�c�S���ah�$eц��ƔP'%-C�b��nw���9;�/�)H(sR^92��C�r�"��v�/�u�v֎�|��5��G^�$ � 0�	�,+,�61��NI������O���]�F��*-��Oa34�ж��'��|�U��{��E
~Al��t+���ʻ�!⮸?��$�i�F����A-�?[���Bn�KK-��o��'fXOU�� �C�t��
y1PdM���87��+�xPp�uizk����cYf�MMr�/�A��pbw�+m���֮����U%��H�8��<���ǁ�fY���y7����J}�n��������$}b� mX��n��2ӳ]�!��V�D���Xb6e]��|#9�K*�˸�ƪ�K2�
�H)�ĂPysyn���A�I�׷�՛�kļh� %G���&��SL?Bo�G�\�Uy�'�E-�<��{�ϟS�q_�ܧ$ǧ��Fl�Zu����$ﺭ*7sxY�E��S鎲���EV\AG��FaS�y�w�1�ǯ7��6�9�HOOM�(�Ȉ�_;~#ppp��Ͱ~o��Bh[�R�"�p��c_\Z�{��i�����?
�d�\7����A�:�����mT�������K��:{����=���-�>���;g1�4@�G��3�a9S�<[ ns�1���V������ߺ�]���ibē��2(Omp�)R��w8s�w�˘�b9}J�R��m���ۻv��&�uƹw�'����x������!�un�[	ɏ�����p�ٶ;c����M��s���Оm'Fd}��>?S`T�\�)#>ƙ��,�������*�,Ժ9ί��{s4*4A$^�Ò`a|.U1�ں	%Q�����iF����ž Nᆲ%_�[��=�n�!��K$444�ᅇ������~g|�mil@�|�m��$�2�l��1c?4��yh�u�0?-��υRn�[�{�2���~�̒�f���iFK� �'��nZ#��$��}�2z��w�'
�����������k��/�QY�_�FFFp ��Tmu|?�����r������j����, Q$��ߚ��1-�yOD�;��Uң��-+)�5|����H���Dr���q�aA��� kBd�
�l�lI�=L��i�t��K�/�Q���W�.��e���a-��u03�.	A��s?�4{�3Ʈ�p��yUbA'�ڡ�Hz�\,;ŏ��>�~�e�=ߍU���DLUS�b8B�)���S�������l�P�v��1�rݱ���+�7�0�ÿ�a�=?
̉t�>�ZK�|[����|�ٔ�R_���;�n��i`іt~���t���8��i��jMo���qJs(���o�՜����Z�U1�4K��Vv�R��}���Q����y'b=�8T*�M'B��(������<�,Hd:��M�R[�%Avo��xP��S�G?��u&�]��̣~�����t�z��㩐�
�HmZ���->vC�g�hE�Z	�݄���y���n���� �9�����S��ەu�ϖ#�p�����/!K:C�mSSSMp� [���(Ԙ���j6��w^lO��j.�J�g�An�_Y��{��|�_�i�C(�1�FM��]�1&GF�c�袸d|;��)0D'6�?����gIv؛�E� �0����{���놾� �_���C��6��V5�/����,2�}�vs޷�?Y� i���-٫�>>�]@�7o�_ERWV�#v�����|[��{�! 넅�O��?�Eka�G�*�k�9�Њ�/����R��Y�΅����J��hQ��M,k2�k�骋×?�NW{z?�O912bK��P�n#�aogBW
x^˞��:�_l���BnsU��U����0O���T�V$e� 2�_�O�+�ׅ�� J NV���l�e��ֻP���ɉq&3�s�s]/�o#P����ĉ��!m��=^��@ux�{iݰ�Rٖz���������,/:tn˭=���:$�G���c�%9!�U��NU�( n��s�zD~̢v��r�W��~=|���I�7�Ym�=��r��uA�ybי�����%1Q�AA`:���oT!,��T��Er�0N� ��?�-�-��߲��GVWW�B�o��Yj���k=[2��n8h�w��hPQ~lm���9��tB��8U��J��>�K�ݺ�4����?����_KoH��Q�q*�pdR������d���4��4�����-��ӧ�x;����<�x ��g����vvM��/^cy���׊0���+k\1�F�ūO$̫�d�yä<�yv�j��א)G�O��֝�&���\[<���_��>Da��w͘�iud�%�i.�{=�Z��m	�=IWK�O�WFf!N`9�}��GT���P|ZQ��d�O��#��,,,Me���ӵ��-��0�
�;2�ω�m ��a�v������@��z��x�$�R�W���sx��,�t��*�V���|��� �P/�]Y��y5	�R�JLG�oⲮ�Yu�q�ej�{�����5&�%Y���:l�#����*7��9�=dM-��E~X�)	1��k�[ny� 	9�|�j,.:�2�gF!/�>���u6�L�{���gM��n�i�Z���(t���ް+P$�O��z�؏��b0^uv]f�KgM��ˉY��N��ޯzv�+.�%˕���o�!��U9˒Ѕ��03�) O�0����*Ҡ!��X�*��ϼ�"M!kؿkn�%�=.����I��'P�(�|�����@e�>������p(�i<̫VdG���D��-�OX��}Wi�g�(�����H��q����)kR�3�(�c�(Ae����3n:	�+�;��S�:b���{����޻R=�r|�ժٽ#r ��U���\�R��{���)D��7��5���� �+ �{�8�[����}�R5�u�)\+휃���q�R����c�l�B��w�;�o��Չ�B���̚dr�����{�֔O�t2�Uf��Y�r�Ui�kQSoe�&]�Q��²�fE,N*�<�]��瓅�-��o�E�O#s]�	.�c�?�'*?�����p_8�rZ*s�wlm�Y�S�26�Dn7���n������q��@��Y�5?�Y*����n����h��5Z_�ʦR���x�}���0��t�WXk�"���_�`6�0��@������6vH��x�:
����WȞ�+��t/q%c�e��E���n�BG��(�ރ�o�[�dY#�*6�Gb(V���[�g�;�s$ԉVbW}^F����Xtj�����pI,u�����,���P� B�� �k��J�R��H#���bP��8��@�d��˞{�?�C���F�NoD/u{f�T9�eI�c_�:�������{<Rf̨v�]�X��	��_�w�+m*.-}V��cL���Й���)�����q�9��(|�ԅ���D2Z���:.��Y��I*]��˰�N6p9�Y�t`�P����W����o�5�N8E���¬+?�!y���+j#h�q���691ͪ!8߲��	��]sb��T��5�.E�ݑ���b�BӽJjz�w�(�I��}��GNP�!Y���*	��a��0H �|���ъa��`�l���?��J�y��mhk��'6k�o�k�����yW��� ���9|�j�C��d>gQ=ZWf��@�q�O�������'���#�1nQ��w��{�ݚ��|b�W�驽F7Z�W���o�!M�,��+ W}�]G��|�g�_^EI��Os���+[$V��N���b�y9�YS��]����m{�UdHwh��A{gu�.��\hf�C�,����}|�<��=:S��=���J���)�i�Qf�6\Sw���gXJz&[#smOF�0�|��7�q��u��d�e/ŚB�Ӎ�O�)��h�,H��Y�[��94J�>�9$�*݋Hs6V5�NcʫA:T&"���b���<�B�+%�Q���c�>��ޑ����0x�.0 *U55�哈���gc��d�"��@��Ch��!6
`5jF�P��=��R��i�Y�=�<�OP�ɪ�v��{���zc�돗C&��&G������^1��gХ��i�"�� P��2����4�+P���Q�����HK����E(C�R�.�DK��F����v�r�®۩���t��+"�9�Z��H�.�z�VGޅ��DNL0�W">Y�L����1����᫟����U0Q YXs� �j��W��y�V�밶������X@@���tWH6��	q�(�Ql"5ڃ:�SV�!��{��#����_�7�2�q��zWű�9�*�$��Y�q P����z�,��Q�4�r���|�5̹�M%�XMuh��au�E*��U���<x���(�[���vq���ԳN/���$��k)�?ӧ����@ ��LC�P�a������]�������{�Ph:Yd+�v����e�Kˋ��m��7����
�2y�8��7�<���,k�:�W�]R�D�y�]�ؑ��'�=��7h�M��g��r���τ��!����ޗ�Cپ�ߖ"���,E�-�mdW�I�BȾ3�,m�]��K���}�RȾdF�d�����n�������{��q<�������y]�u���u���N%������f��E�a��4qk�W�-_�!b^���۰(���f�����ូk�f��Not��	ujpHjqgVxsq�>� ����?<��BI�I!s�ک�{o��<�5��me�<aS����X�v���mК�暪*�ʻ���7-�ur��/F����?zfÖ�O%��)�[��B0m�J�����8�ݍ��=��O�b5^>�g���ə���c�$;{!'&�ܾ���]?M�5��������.�٤�c ^�$�Kn(׺Sݞ6���y�Z8~z���C�}��śO�	���S�s�VA����w�D5��T�>����x`���z^�\I�3Dڨ�����Ck6��8��$Ѥ��E�t9�ڰ�,_���o��T�K���Q�γRZ�9�m^*�'���iB�n0m5�ul���$c��*%�I�ۡ�g#mr*�����~l���5{��΢��K*ö~��u_	;&��3�b�qC?T��|/K��k}c@�6m�IF��N׳<���QW��^� ������a�V�1DO�S<1�Ǘ����f�B<p0�ݠo��j�Z�<v�	�!Z3%e8*��+�∵�X����<�0%�����Ԛ)"}(�
�Ic�7�9�g������L:Z~.��yV�մ=T�J�Z�y�N.��!�f����Z^y$v1�Ԯ��a+����9��h�
H|ll�rn��Y��)��@W�W"s�h!y�S���m�-s½�/����/�n��_�қ^�!:��(,5��-ќy��YkR�9�g%�:�WOl˃��B���}w��ꐅu��Y��`�qr��8}��
h�]f��}� �'��L�j�I'�ʑ�9}lY��rq��x:ؖ�_>���]Q�E0b0 ^6ӧ�mWc|���R��
��|����{+a?G|%�f��㽁���E�A�Iei�5M|���$p��]ro���UI���vЋ��5~���Y4;;9�ORhGU���y�OҚA�+������}��9�{|ksSSS�tC'�Q I1{�y	aښ/��[e�u	4�hA`�Z�o�b���ܼ����9^��T�N�2x��ě���L�e8���G�7�.|km  B|�Ln�������m4�"?���|U}a���:��e6�������y8u�~g����c���wnBk�wץZ��8�}1�B߫a�U��ԭ�Ǖ��˓��|k�|eH�Eݍo�+6le�Ga4^�+��@�(y;/�S>L�ti`���b�f7�'�TR83�\����"�����;�I���f�:\��hSa�*69���.D�3~���n��j�7��}%H�Fr)A�Oȏ�����5�~�i_0'�����v��(��n�\��o�7��ˢ�7`�
���δѥ�}�)���AZ�������ܨ_p0D l�Z��������P;�D�ci��v��:&������G��de����/��[~��<��mT�����(`�x$bl�'�VY�]PUE1_�(�)��0m�ɴa[x��4��o��r��蜱���B͙�pY���Tߕ�^��S��W�"�����>�]P�۰ck�Y/ؙ�&�Yi�&A2�׾�:�QS��?.���Qh���ߥ���iK.�����s+U���}��=#j��rS��1��e�ɻd���<*gA3�^��?�	��~g�ڨ���r{Q��IT}�����o��.o��X�b���׹����2f���N��N���~�aj���SK�>;/���u���)Rlѧ���Ŧp�͈�*�D��˶ʅ/��*�>���2L����9�L�6}���>���%��ϥ �ȟ;M�'���������_S-�i��Ub��O�ڔM�ˊFG̸���?����0���*�R���;�<�Q<N[��^���+�&���h)1�}�%ɧF��xg�O�W�_�W�����ž:ޯ�c{!��
�_^�v��X޷���9 м��Hw]W��`�ō�^a�grC��P�J��ݐK%�@t'xrl�,��+gY��&W1�uQ�H���l�o�p	k?��U��
��ak�~�JTD�g�T?���$&}�����n��<m���_E�Q�&�e�|*��5������$�<���R`L'ڙ-}n������h�*���4ԥ�@<)%e	d�a�1U�Isx�h�#X'۰�1�"���9?�u��Z�ЪU]�ᅕ]*�R�uZx�x�ҙ*6y���;ɫ�Z=M�u��Nط?�0�т�4L}I��is���<<�<fD�Z�$�d�����}I
�e1>*�<���J��b���L2�y����d}uF�~�*����b;�oI�07	<�a���z��u
��g�������CBv/��5CY�8�3����8oC�y����Z�6+�ǖ>ΣT�S�s�W�vli� 5y������iw��,��i\�y%������H-���@���[`[���҈uZ��ħ9��-����Z^[[�!B/�J�((%�N��M�C�bT�<Q"��Z��n�"10@n~s�
���TH���F(p)N����w�9G$�;k����o �/��E7���fN�u�-�wL@��hE�:?��l�*6�\�������>�d��L[ ��F�}�H��?�R�`G}��I&J$�a�ϛ�vL#�ܛ���+�Bi�|�A����X�|]]��h�+����A��0"���y�?N�zK�묓��#��y��(ͫ[��ް�3<rM���kc/j��u�P�p��E�N9,_�n��o���`�xy���.zvp$$��%Y�/�4�"�l��1_���`�'���+�ƅC��k������}�,��KO|B��5r���.8�܇k��N1��� ����0F�b�3�Ӧ
�d���B:gs�����qW�O���V�z{Y�V�t&���S�v	O&�6�_�ˁHD�=�mH�7��\4�p����ۊ�#^�8m���.TTTɶz�N�w��Oz����,umr�p@9�w�>��qd$������Q!�:�m7��9-������π�6M	�>=Id�n�ܗ��Dh1����V��D��&M��9\`q�n��ƛ2A`s�6�0���CY��m1�25;E�pw4���5�s'�b.�N9���� �{��@s��MeS;�P%��~��I�o�z�U�-�� I��@|,{�"4�w���>5Q����T~��Ʌ�W�c��Uk�T�������^񔧟N��:M�x�;�zW"�YI�/sxʍo˩�G�gھv8��L��.�_�$�h��Z�L��i�(\��s��(���j!By:�WQ2��eE�0$A���v�Ӄ��x�HQp�Aٖ��0|6�X�o|��h�lw�Eq4Y�,����u�������I���Y��f�ZUz�,�a!~�� H�o�gn��W��uy�_��lo�Ē��G��[W���"�pn�����#�m��x"�oR(uȲ�,t<kp!�/h�^c�eᑡ����clI�'�%�_+�|������G�Bw�ϓk^F�jR�^6�w^I�H�\C)���%STZ���L�3�~R��*A��o�3��U(I���Q2�� 9Z6� ̈́\6o	>�4�o�p��Z��GXwO+\��j|!���
�8z;v^���1��0����h�h�FӪ�9v�o	����#U�z�� s�	� =�R�V}�~���i#����Z��(���SR�U� :�]�H�P<L�%�Ѫp ��+����/U����ӿ�%8��x��VD�Rcf:,�7�A��D���/�C#&�m��*w�=�^�^����B6W���9_�����X� �*;��٨Xu(�y?��E̻֫�&�����������P:+�O�t ��$H�[����P�t-�kY�8��4����Oi!�׾q2izi��T�����0�N*(�ˎޭm�����/_��������)���sp�˴��k���.@;�ҕp��m�$Y�0�F���TZ�����y[nց�H9Z'V�«B����-�}�3]��K�(> �⤤$�[�P���*;��Fir��7K���1#|KM�@ ���"�����v�@`��};�T��F�`�J����lDۓ
��b��pW(�����b�jy�7�O��k�S���}�7W�sIu��ґ�(����7D���s�����,*1���W-���2��M�/8���X�	F�Db����ȳ��<�K��.� b�f�� �����Y�g�o�Q���1�h}>] �'|�!ܚ�֕W�	�ݝ$����8��M��v~����;�V�n��w�[�L���Y�`�d�חJ�X�Q#厽��&�Q�N�ir�ip�9q�7Q�1��t��β�$�6�q��|"�L��t���g���T=1��"�����}&|N!�����d�,�S� �k�6��Hq69%ٱ�A�đV��qp,Ҵke�Ѓ$9p�vA8�v�����c]*9�����H�k�&���/����B���`2|{U6�/�z]O��p��5/B�'����6<<<-�L�::">�X�y��(�>-���y�OjZ����^���J �����`g�0㶧?LS�)��b�giii� �Y��?'��F	CV��� �(�O�^K�^&�	�|mȃ]2cp�f��0Y[�؏a��"�W
�#��Hs=�|�����{�^*I?�S9�
��ڇ襣� s{�Z�n�V'�����'�B]q���o�������75�ɶ�'��8��#&R�n2 T]M�:d���[�m�!a�s��%�b�\�@�<�I��������73`&�����P(�a@������Lx�����؇3˼��U�k�Z���`J��#����+`�y��ڟ���v���a@�]��;g��@a��i}9���4��6oU���¡��N���`�n��3#f�������� ҿ��X;��W^^.lw��(��BO#,?�A�^�z")ēW�Z�� }��d�<�-ť�J�*�?/賘LX�^b;�7���6c����(�g��Ļr�*)����<�
�G�V�P8��I�b��,��O#� �ңv��@���[FF�0�#(W��rP��g���WO%�W�����[�4�d)6m�������J�A�J�U���⩩)��z��G/���[�$c�}w�F�=��=��ś�WXlV�33�^�b�9��,���ױ2q27�=�P�s�𢬬�r�D�&�T�9���/b�U��4����Q�X�>�ꙣ sF�6m�|՟����f��������Fʿ5@��ЁE%���Ha��5�yg�\��`��.6y���1�^�1�T����%�ȪԱ7KǵrD�Z+[�Y L����`��X��&j���u�G6`�1 ���lF�9���0��uD�w&�Ԣ�z�@��j�tz����%{� q肨U�<:Ќp���{R�J1$��nO"�l��Q�a�p����μ�}�J�T�ej�z2�=�A�k�{"��B�sh�f�x0�w����ol�7kÕ�Ús�}p0rMa��أL����v;f ��"�
��|}}�oP�����?χbV-�R�ܨU�u�Ȁ�zt���"s�|��k� �~�Z3�r��n�'S�W7W�ws>'�1(+��9-i27Z��8`u���w�`r�b�@RR T\�ܙ���|;=,	�������o���i���̺�=��<"�&�l�;C�ȧ"�]A��ٰu�p����bm=��XQY.*�y�fJ����"PZʿ��a�{�����c�.{�	��~���~*r��>&���ӧ����=�^�%c�㙑�Q/��؎r��e��#s�hq;�E����WO�yӂ5n�M{+������U�
��3���Ӛ6�4�FG[{�0W g�d߽7�ܣU���|J��A��Y�5.���DO+����k~vI�×Ce$���^j6�临�^�>������h
�g��ۨ_'�(�E0t��(����ĵ�#꼳>��`�Ys��7)��H����AR1�W�{�EY�����*) ���Y���v��K�w���1��;2A������+�)r-�NW�Wt�==@ l�>���x� j�:�X��)�fQ�۷y�������fV��=��)�bmy`��p�l��7��B���� �R.�c�q��5gA��I��x��-�8
=�f�JX��E��W�DϦ�0k9��s"������R:<5D�xz��ꐟ��ڢX��T��c�֗8�Rw������jǄ�Ba���F����ԌKġ$m���]��P�����β|vp��m侩��	R��[#�C���0˯��� {���'
����'a(���Bɿ�|;�ٹѪI7s�EK G�9��\M9�X�'�_M�1�)��`����D��{�� 2�Y�\�L�PX0~�!�-qZ8�F�yR��x]j��Q��!Ҁ-RZN�k1Ț��s���ʔ?��)3h�e�%!n��K�1������3^�|���ر�ҕGj��nWŻ����*��i��Y�2�3�v�"J���.X j�Ȼ���G��{���������dU�Q�O�*���,K�����ٮ���-�r�x�u8����w�ނ������g�v��H�>J�7N���1Ɩ��Ο$��6�������j/ʀt]��<;5&爝�]�h�N�n�ۜ�ԯ�ԓ�,7�lߙ�����ÅZ`����6.Z�ꖸ�*���G�� �)m�~Y�l�����+����������՗�=��ٙ���r� X��3�-�i+�*>�
����r���d,����^s$҃-AЦ����b�e�Ww�UT2/݀?����$��p�R�E�.t���)�c��\�G��-&3��C|3JEL�N�����i���J����t%��@W8�q�D�β	�PN��tuE���=:��h�j��J%����XH��6	L[�xiEEa� a0�(����E�����2�2U����A_��������1�mil�=�ב�/�[y�h|D�����O�oV�,�H���n`�e u����*%[@�V{N�<�L����x�ߟ!�C��G˝����Ƣ���Ē�WF*I��JIF��r�;��{�
���u�R@��9XQ8ο�7����)x�T��yT�>v���I�%gi���4���`�x��Y�[d.��ZOp^TN��͝͡rW�e�	�pt��g���-��P_1Dn8���Ӝ�e�|�����.���7�c��tL�-��#�A���-ߟ����Q0zn��S#�Q��c����
	��;{V�fxg��}�Gb�}��͡Z>��U�Slo>��@$%(�׮ ʖoo��L<�×u -'��E��P|�Fь,5�{B u��5��pttĚ
Z��F�`���h'G������o$p�%b�.��/��'��L�?��$`xt��F��!�n�끮����'{
�� MҘ������? (إ�˂7\JEE��OC�B�[��n~/�;���9�P��g]8d��X��Hџk���I2��o�c�;[-	*5����6���Ey�M�6o������<<�X0)��]�R�>�����xv�)��I�h�'�����t������j��Gih�P�P�91߹S���ԈBL��4>?2�{/���G' )��a["s������׋���O�ܻ�x�BJh@:%�wx_ �_�@��"N/I?>9�V���i��+�tZ[[�em�z�y���]]W>ݠ�"��^�L�����$�7�v�yJ�*���LД�J��Y5�;;;ؒ������Rz��|	����+��E���Y����������B��<�0���H)((�V����{� ����w_�b��1�"��K���_ ��]*Ӯ�r�֭�_}	�/H�{ҵ��� w3�f,�)ia��`�E�Dz�E!�������TʱTj^L߽������߿�p�i�g��6������1� X�u��衲"�6oCТ�����Sp�j��OI�����-W�gϞ��� ���ݐ����RFz��3��K/�
�<t��c���S��%!$��W=gY�T`�6)!�9�#I?	2k�	�N��S�Ⱦ��::���5fsl�[ �.������/���sIu�85 �~��I����d������<�|�4�-���Eރ-���}��oe�{�5Q4Ȯ��y,�q��q��O���+-Fzf��a��������e7@���4m��6�3�_O%Jt���Z�����b�����U��msh�!�����%>������020 !y�\���+_+Q����N��@�5� �)��B��y���'�|| ��l��=���R7�%~�J6.�w�j7l��t�P`J]*�lUf�ł l;���&+�>���2z�g��y���/O����ZH�2����O$���_�dccK�-}a��ֱ!���,���/�ډ�>��Ă`��,^;�9�,x�ω8�ZQ0w���i���V�|U򉐛G=gG �G� s��/_:o�& 
���]_<������d�ȣK6�"��?3C!ȫ(��YY� �1 �i��WP����� bU>�?�َ���e< ���ԕk�,��qq����z&'fy�t�@���'���V[�tq%�{W�J��׼�n��_X�Mvn�L�����#���*�z�933�e9�RW�����2h��h�8t�*�l�E�c ���ڰ����R�^Т�bk̗��=�&���r�
��P\$�jh�<���-�}mR�w�Zl���� W���\���q��H�� ]����H�����zl�E�i��L���?��L�M�m��@��Y=_؆fX�՟[/(�t��DڼNlr����"��Y��7PA���^����C.~�7%�5X�$���lP�˃��o\���횽��� �ET!�1 ���S}��BBc��%��e�z�ak5`�|�̷(��<I��w0����lU�+��r�c�w��%�g�&?w���"�677�o^Hiz��	�%D0��\�h\'�n�xw2�?������cg�Y�C�b�?�N�d�3#���5��. U��珬u;�<4�*F<�	�x~#8�k������Ǐ�H�h�U(�ʻHx�2�)���ܼ0��*����ΛUnA
J$��T�Tֹ�Z9���X6fb8�X*�7�Qg��5a\lbok{��S��PsSy�����}���5��K;��}�SQh�o��@�!BU�fȧt��V��v��X�!�]BѼ���a�-�a�9�����y�sO���U�,�x|�m���>�;��Ɛi�C�W��֍��I@1����w�9Vi�)q���,I˞�;����;�~�x���.�TWrFAW;���Ms�T�|7�|s��~��ma�������ߠ��&T�Dn4bC�#?ց���6�F�W�� I��XK>�s�r�+�#IT�k/ī�J�H��SAHm2Ѥ�{(�Gk�r@�����
O�;��:�w�|f�����`c�`�2i�+��t��bqv�>N�0U�Yp�!Kbrӈ9	�m�ƨ���U)z�VL{�}b{�.Q�}Q��́���سx}��=+��.�������3��x]���7�$r�;��P�7(�+J M�p^�7��b�"��B�Eҷ.��{�~��C_���1=oj�ȳN�7�v6��6ofN�WD�{�o��,Yd��k���U�+�{N޼!Z;�vÃ_qW����_6ȷ��>{� � �.=�@]�tm��G�t."�q�틁C�H�(|���M����ϳ�1N&
�@��VN�~�]�������ԕ���r����PČ {�Bp�Q�����{P��
t��9��L��鐫SB!�ӧ��k5��q�L=�筡'i�o2�>��4�d,��m"�U��n�`�'%<��E,�M�;H����ǚ�Sk�е�d&ocW����d[w$�[&�B�s����S�+4�q�>��s��P�6bf��-�o߉M�l%b+����+2���7"���y��,eA�O^�x�pR�ٿھC	���wnv bB!Ӌ���?��4�f�-��$IIa7��ڎBfW�z�<�j����1��&U�4P[N�!�nHjG�l�s�&��!�@'�䢿S��ڮ`��f���tYg
�X�=���47̕�H����6�K������!g�Rj��Se\�Z0隷��VVw��B>jU��u�G�m���b�w�M�)~�u's�2ᭀO��uTgJ6�.�h�R�R�1����|i%���7Mb aop&������Y+�P��#�U��m�-��v.�H�5�)����c��'��!^�nº�5�v�JEHm=[$�}±���3t����"��������ϲ�AN�3�s|���4i7j^5Pq>ZO���&Z.2�;e�J&K�n�O�^��)m��b��Q|��Ӓ�=��?�^���/����$��eñ;�"�z7�\x��� P7>?%�v���^�@>&%xe��;��pJTs�
\��������ǜ_�y{a!�v{X�D>\�<���QI�~�-F(1S6��4S�%���}�h��DF�K�!@��Ȟ��k��-��[��v�����=�*5����VEA������h��[�v�O'���+9��v�aD	���h�Qea�U��*�Ͱ!���/��`z��:73���=_q���*�����M�.��x\$G��\��%)�у����V�{�V�^�˙9�W}�p��Oa[V^eɕ�)r,as�Z��+����x;t�6p%		��׶_?6��f�r�T0�r�:��o�P�Y/�V���3�sۘ�HH�9�+��Lo���M���;T(pF���E����"3n$)v�!��^m��]g��J�Ir�y#'��!T�Txy�t��sy���9���w�K����e��o�}T>���h�8z_��#B�__ʥk���+���������z�7[�*M��k�.-M�oTk�/�O+@�@k�v;���FIDN���Eƕ�����:�@;y�Qo��pv���'��M�]��Ic
�ߑ&���x�rFL<��t��8NhG|<vő�O^�ͫ��HhW����B>�$��/?�:%�K%�?�D���4���|���`�ؼ���E����3!�g�R�:Ӑ[rEhZ�͖�1�M�i����D���/LP����������~�L�o�w�,9}|_�!�Nuc�!���:jO}
��'�=rW�h�%+A3�h}������O��\�w�
��U��#��PEDQo���.��NS�,X��.,wO����ڂ�Q  ��c�[��t���V��mo�O�4�S���3�Go��0�tQ@1�9T���Kx<'����f4����'}R4B f��7��e�x^�=�X��י����?�G�{�� ��f[)b�B�y������`Kc�v�(hM��w�O�i�"P\�i��H�!�{����_q>� Z�� ��'ϨE;%
 �U�v����Xq�z�~vg�T���w1ֳ/�P����9_�Z����&m��3�>k+��$4�?a�!��rN�$����N��z:�6���9B��In�e�i�L楝�hT�Iq�������ν"�c/��2]®zZ��C��h�:?�.���t1��w�rY�-i#v�r��c��f��=\�˾ɮ�C� ��v��7?N/�IM�<�C!
���i��3-�F�0��o���v�2�Ҵ${����0��̇���R�]lL3?0�����Kv�:j�
�>
̿���.,��b��E�B��i�v^��T<��DJ跚�t�zwψ֙�9B��X���L�o}њu�.3G>�H��Z�9k�G�u�M����ؖV�����T�r�+G/ϩ�:�Ϻ��XD��T�Q��d��y�p�T ��ں���~�sx�je�}�$ў�B����`�Bu��-.�z67P�1ዩ@��&޿���6�T�&f�9\�maLr,�٫aF�4�Z<h�G��F%t~����9�L�rS�,��cK���:G9��F޼z|(i��Rח������BK�YdfLD>�ɐ�^�1�6ƛA��
���VY����CB�L��*�����u��?���_U��y�c�\���δ���i����_�O�2���ޥ�oP]��G1^o�u��>f�!�S�o��@[���ě��*�6eV�_�����.*+��Z��Mb���7ʾ~څL�0T{';���[���>�	�����h��g���f��r���:��ʙl�t����5B�<���9�t�o��l�Doɘ����,��8Q��ax�Yc�����r&�>�߶�'u�z�[x�$��#��*AD���M+���	VR�L��p�Ж��E��B��ʀ��y879���щ*,75F���L%o}��X�o��WAv����7KT��:��ݑ�Lo�3��0ŏ
��"�6�G��E*K\�=��+<l��P��1~���͜J�k��j�^�>T?l�Y������i�Կq� ���yHZ�|c�����*��{������*�]�(���Ьbe�=��,U�:��|ྴ��*�|'�o/���Z���N<������K�>K�k��gI�!,�Hd��ʫ��7M_oL���Io�(�	��S�sj���7]x���. �Jzk��Be���e8�-�^��O���ȩ8�NO�g�?�$2����6���O}�3�\����n|��]�_��G��{�i��x����KKW'BY�CN�R@㑀j��;j$v���2�<��`
�)�d�	��K�����9�_sm�pF0
�P��,	r�M�]�p�+Z`b�_��d�걦�l�7��n0_:�u������V�Gb��^,��ty{.�
J��u$�B9�l���?��Հ���7���×��F�1�O|"��k�<�p���S��o���P(�����6������&���!h퇩4�����Qh�����j?l��k���w,�������/7��p-N�Ev^� ˕�����?
����}�,A�:���=���dA��Jƾ��@+/����p�ߵx<���B����?}��}�*������o]�����g"O��"���|��@�O�N�d�TQ(��&�����Io�ǹs H���[���կe�Ћ�_򑑑.|k(���X��!��縡��*��^�Gr��D,fh���mM�D�@}����WX:�J��!��phM��)�E��'}�������[u��0���=$s���]\l��"�obuĲ"���A�k�Z��Y_m,w'X��(�A����*�q�@���.x�T��l��+�����(�tJL"� ���[��A�<T�*���g��8,_a��("��pԖ��ќL�0�R�p!)�j�*���{�^��;(��u�"Q���:��&h��mN�cZ�&�~[~1��^ú3����1�����ګ@���ˊ�1�V���_��Df�D{=(���꽆	������������w�C ��̓��Z��g�ӗ�K�h�>�;j�2��z�;�uS7�� }3x�'TD-n����ɬ��^�|
A�A|lC҅��YuG�3��>�1c�xJဗo�=l�a�b�[3&(�r�ۯ�m����SO�C�����u~M�;y|>�����c:w����DSc��_�]J�1%}E�J�z���20�$�4�ɮ���>��j���Hg.��8U$y�;:P3��H���8���i�_��J'p��dp�Ӟx�M�\���ЫY�RE(��z�m瑕e�/�M,4È$�j�{Q��"����(dV�z+`\'�=I{��Ƴ����2bWj�H������K#��7%7��=�
�W ��
���ۓx�p}ͮ9bؘ����l�&v (�������\���g�=�~�(�����:d�A�@"�=	�e��y"���n�B���N,)K���G�;���	%h?
�-�r���z�@p4�Y��H��8��v&�<�(���U���O�`�ڧɺ����,�K�oG�b@�N��g�=]w�$oGD���W�><��+2;�cͱ����F[�H:�������w���C�½f�Ǐ�7ҡ>axj������"�Z��c�7�OjF�و�>f���dgw�k|�3�ξyq&(�Z�`q��)q��'��xE����
� �ѓ��g���k�����\���{��������߃�.\�}����m���L#G���?��"4OfR�k�b�l,��������}n<&#��lN�yTy��ҵ*�ң�I}�jZ�{i�d��p2d������ǮU�D��3��-�w,��Ê�6��4DY�_�^��g>w��NV��)I�J>.�r���B���ndP�mp'�똱�0&�w� �6��uz�|o����1d���oOY�OH�m�I�����f.�C��T����	��ËJV'�='OO�3�0>�w�M2O�4�cBJ�s1�A-�r�Wl�c�}Pv�m��k�^e'�2+�/���r��seO����X�f7�?nm1Ⱥ���W�͌&2� !�PP��6������q��\m&ˉ$ ���O:�C�f�4W�z����w�j����zk���F32�� U���\�֏AY�iozf��7\7��W�L�zE���~dȇ/?���1�� n����f�L,�5O�h#���e�?=ӻ�������潻��R��USY��WL�v��+bf�7�v�TM���g'L��׆�f�����\�����k�����ݕ���R����$ܐO�½��bT�f#�{p����4%5�_��5���_��5���_��5���_��5��li����~��{��D��@Pp<�����c�Ǯ�ɷm`��&.Է?4�'3����V�4sU$�HW\�����xgg��L��~��ge���A录���nQ���_ʩA��}
e��`��l�t�������vh��f��B��V�AF��c��Z��L�!m����w�s�)dV�^�彏o&���g�~�3T�_hOJ�|9{�inߵd�k����YJ'����tj˸vv&x�iCY F^�����y��ڹ4,qe"d�''1de�RX�P=��%�]��� �F��V6#k��Ǧ��3ʭ������
{y�2�ۛ*7J��.7��x�"o������\L�j[\$����)��d&��Lh<^�k��Z\\�n�{�h���ǱZD��5���`������{P��XH��ٴ�~"���4.i0x�.v��e&qke�n�C�MZ~9{q��th׹qY����=�>�$��vNkRn��K��EH +B�򃲌��?-�W2�h�O�P��4�P�x���ij�.ݾ� PK   �rZ$�8�l  �  /   images/aa130aff-16e6-4627-9689-819d55b5861f.png�YUL
��Xq-EY܊����K���a�RtY�_����;��kq}����M2s�9�L2�3�/Z��X�XHHH��Jr�h��[0��Ÿxl���d������?�m����p���d��e�j�����e������ي���&�D�	�F_YN����3�z����k����Ԏ����(�Gǳ��R��7���c�JMNf������a�\w��{�I���kD�b�K@�)u+h��,?I9=̚;�����[�(6-�r�d��CGG�%��+��1A������G �����B���	�A�eF,M��Lo���k�=�8%_<�3��5���K4�AlaA��~��V����6�~nU���٤�:Ƌ]��d*
����W��CMy(%.KL�)�U~3"`��&���Y�t t�I� �Be���qkP��r�<f|0$L(��-+_�a�� m���$�J&�a���%���}$?�}}����4��ۏ��˜
|<gX��m�/���&�f27��+F�lȏf�{L�4d
�"��)"eN��_���`��N� �W��ܥ��d
ڵ��Ϳ:��-�^���X*�^�☈"G��oւ��^���i2���n	�ii��}I� ��M�L_�n
k|��g�^�D���Fg�Y�U��'�Ԥ��������$k_{���A��G�1�F\���uGLvaf��<V��W��f^���2=Wt���\C<�m&�	@�Z�O���g4��͆R����թ�#�7�Ȇ�A&��f�vf5
�"����0��hż_�z�@o*���I�3Mu�l#�c
���H�Z�I�C3n���6���ﴪ�	�,�@_�7���E_��~��ܫ�[&�N4�X��������'I��^��D��;�d C�uI'��;�����L��ږ��!�@7�<�^�����	�ʉ��!Zv�pt6�L(�QbG���Y��XHZ�e�<Z�L�$��K�V�jN]��{��i[E3<ӿ����R¼�`�ӡs@^��pv�Z�#�A��4d!~�D��޳%�{����i)�*7�CՐ��\,��{�_{A���>�Mu]hm�w�bD!�$_`�12Ő�Y�D	�,��&���W;��uo��oX���N��������c����`j������{���c�sH8�0'ޠ<C�ȲL�Q�ۗy�ߡ`��#��Q� ��y��IX��L�J�{�X3�̓0�1�|'��f�9�CC�U{�'T�K�c0�W�&O�BMJ�7&�꠰l�j��������X.7��k���leY#zu9`�4;��w�}U�@�l�`V�[�Zl|D`�eJm�c嶚��lnQ|l��;�l-��|�8�Z�-b�P˪W3��OIƭq�:��KS��d�iؤ�)��)hDסQ����UU��e�K��iKR��@�^9���� ���7G��*�p6�����Ir����1�q3��	
�Fl�I�=m�h	� }9!��m�W�:�1�jC�����w�(��b�������l7��2�~xJ�֛}���F\��w.5��ߔ�h)UV|il��;��cL�{K��ty��{ �``���C��p�w�kz�����I��g�'y�h=;�@�D�{:j^.�m⅊��|Ǚ9����;R�ȍ�� 3����xw\���CTl�y�,u�v�e����Y�(Tc4@X�l?��%:��v�M�(��� 8�TZ6�[��_��Rz�#�E)��i�{�5��.�X�uj}\m�w��~&�e/���H�8���Q�/���H�R��5���_�5�q��i�V��;���~�++�9Q����9=�CK�;G�T�N��㥲b�=;�p��>�3���W��.1���E�����|��Kv4/�t��XTJ��6�u{��%Ǻҟ.���G@���:� ��y%��
��E�N7(�� 2�-���]�H���Z�  O3�*韭�<m\�����t�pz�#�����Ց��Um���C�nĮ�$�e����uesM�����?����pc"a�4u�hi� L���(|�ϯI�L� f'�E"��*٩��ծ� 9�-]�]�������S�;iSKn`Uȏ�=����R��8�b�96K�A�E8�կD�h�⢛ns�/4��b�#5���6�R^&h`�j�y�9w�T��ێ�Gy�x˞�iz
z箹�c�*�_�9��Rg��U]���,.V�m
g�H ��rK[}����цQ�I��X�H�����rZ�y~ 
�6M��
򗢧���A7��!ܡ1�@��I�ĩ`!�j}���%h�	Hm=M��ğ2�2���I	��F��[�!�Myv�LE)v��� 3���>�xj�+�Ҹ��_��a^�h�$�ՖL����q�Rf�.��� ~D��O(h7G#�<qF�[)�������k�mFG7fL�o��k�1ջK����r�W��o���2Q	-��k�z�Phiѕ��"0����u��{���blRxk\�SK�.wFM=gx�)���;��(DCR���=���}���ST�P؜f���M��9M��X��Jlָ�.�1Bf�b�^�����g���H��(�_��_���	�F�(�P��}�y�&(�$՜D�Կ!u�y����e��a��,2�R;���ٯ��=����"3[	���6�rm�E?\L#vO0Q�3g��ˁ��m93X��GS�=]��F7/�=6��z�|�y��0�7�#�����7�}m���4t��`���H�袟���P�N�ɖ��{[���4xʨaO�K3\�qd`��R��sL$����;QE�I��G)o�LQ�uz+v׺,��L��X����%�\��p34p��Ѩ5 �j��Z��g�<6�^ܘ��岓d$^I�@//�!R}�V2qPN��H��b5~�q�@ ��>Jɒ��3��?9��yb�Yř��s���1]%���Pf���&O��O�X�����S���cܹlb��Ya��@E>��7X>�J,#�В��s�*.i�JeyL�P��N���	�@׾q��/"�M�))��u�:�����T؃ZV&���b��(��h5�]�+��9��0�Y`/��|�~�<�����d+�_?{����@�U��bꎘ�״$�P�`oP��R`]���;1�9<P���Ιd��`��rCF"���\ջ�(d>�M%DiJ+(63�Cb|"&��x�xL2%ѼZ����CV(�(�aW`��m��R�E�o�j�SX�r$�h�cz@�S��.������/���kW��z��[���z�K[�tK�f(��z�ôڛ�I�����r��,�*$��;$�|�q���zw���ǜMh =J�"2�Ƥ7���"Q6�˪]p̻�Aզ�s��:�C����w�5�hxa8B�L��n{�?���(�͸nu�$��Lt�z-=
>�EO��M� =�=�pΆ�0٠��Q��e�Q����_����h9>�Q�?O$W�d��/?-��uh�4���)(v�Uh��CJ���/Y+���<�!�Uw�~]PP�����Qǟ:�Ǟu��o0��|j�sv�%�U�d16͉-���Ze��Z�PR�_Y���7�������}���؆X����Q�������)6�	��N*.)>�.�G{��3�L^�u��p)��ÔA�Q��yM����Vp,}(Ll�xh�����---l�PT�ruru�ޥ2c:��n.1�N�\�4�M��3�ť�N,��f�e�����5i�@�Aɭ�-YQ�S���fƎz�
�*w�ÌO�ƪ�����'�J�/���#�%��.���U/��G�+;�ET|VP8�FBM����k�WY"���>ފ�]Rl2�T'�w���QK~���O���҃��b�15fBv���tA��g�q�<QӳRolև̅����A�D�.`7����B���*��R��$�ka]|o[d��J�=Q7�FbnO��I7#b�F���3�|�T�#1��D:��/MV�u��Be������u8T��'�&*�c��/C��̊�|b���,5|%���l�W�d�_���V�{������)���y��4C�dZ s���NX9�[T�W�⍪��ѵ� �"*SPÅ+W!��q#���[Z?��Vl���{�w���	�h�i6�XJ�/��I�\#�)짎��~��x����@�'^�u�! "F}���P�����@f�kM���������`mO��3���((��MƠ5g������본��N��_�b�mjВ��W�O�٩�7W�}I�.N���وa�lF���ʔG���N�$so��]�S�ee���=~뤶��@��N�z�5��:�s���ĕ����R���5֣o���laӗ0���>��^q�������3��2��R�7�$�;;M,ˈ����B�������`��W�p\4�\�qH��� `����1�T)!ؒ�Ak�J��b]��%{���DW$����~ս��F`(��ÑuCg��F�(�+g}}��'��- A��x���6����n���#<�]��a�������{�c��J�,�5�p��qp#��R�ZX�S�/.t�Zr�]A��a�N�(6���_km�mR�c$�<Qq��)~�+���f�Z*pk��Z�f�͞Ff�/eꝻ!Z�@�`ḋ,����?)�*��(�<E"�3/���"���"��o�{�RX�N��/�a��ZU���xm��iX21�:1}�,aS缈M�rwg�xM�u��k�Ѯ��e�k��V���S�Y2�֯�Tw������o���];��nf�/��ŧ�A��\��W�o�@��sފ�H�#��3��m��{"�E�Ӛ�G_�U�]��K�i�,�E���6��tl��$N�J�%9��{�P#6��䓏�#��.�^YSx��WBI���7m��O99.UϹ~!�t������	�[z~� SX]�"{��#���7��4w�M��z���$�o�,lM��u�D�Q���=429~� �����AŚ��Zo�Fc|��a>Bz��
?�.j}�"�F�4�'OdZ-�QB����j�IF���{$��dֵ~�l�EV&y�˩ XXy��DJ��c��_(}��s�T��Ҕ��[��D����Mfod��%������Y��cZ\���$�1�\�Tgp�ڊ��-��I��*p8�C��k��Sm6\�������<� qN�&,&L��0���=��M*�+Nol�X�V�ډ���b΂��z�o�����ӭ�������YĶ��U$��H��)�5�:eW���Z���<��c&j�0�b�m�վ�s���X�O�0!R+"����U%���a��b)�[����z5g��x�$����Ke�����d�@HN����c�܂ח��):__8�$���8�+�Y����JG�짽�4�E�^y��5p\���h��VU٥���h�븏����|��^����ЉO�I5'�V�t=`�},R*G���8Z�]��Bg�X8�F!�E�����t���2;ę����+ݘ�V��L�Cc}����)[�-�� .KfwG���<8^h@`!;��6ͮΒ��z�Z�%݆W�Z>;�[��#���0�%�o~���<;z5D�)a-��X߼}��U����[��̸��W>[��
���D&yY��~�}���cx�3��Ey�1�VC����wv�Ӝ�)1���Ⱦ��L=���V}8�LRo��N� <���5���w��x�4����O�߆��Hc���]H�Z	Qi�{�������ɳG�լٲJ�����̸�V4�$E�2�z�5�|�R�$5R�a�qL�qe��"V������X��	�y_6�IG�41��n����@l"�oz�i�v�ɤ��KlP�*$La��B��g4��i��/��<�:�\]/����d�!`7��k��J�AVf�����Pmܠm�g\|����"݇�P�B�?� �jdԇ�-�#u=
n��m9/.��\����\�]��g5<�����y4�#F��C!;I�@&0S#��T}���wd�@C��{�K�H1��7��,���M/�K>���-N<�6��"�wqN�5���s)��G�q*%���9L�Q��0�wk��w���x>0.A$���-�?�˙6/�PDH���>��2�P����Eiap�13.�U�Yz�C�)|�s�VkV����#(V�ʹK7�������ߗ3S��n��?�p���gҏ8��Bقo�'j���BbZ�%��M;#w�"�⮣c5~���/��IseIu�/�}�m14ƷS��b�#�<��k"Vj�͇�[���V�o묆I��?DoA	�Sv��&��������d�~����6��v��h��=�X�?mΜ��k{�����6�c���W�L}c�w�.�S�~�Y�s�_ٴF�u��;��8���g�����QT�0�ap2�;Z�1''����>���˵X�D�%!�$�ʽc��V�/&^+lB��IJ�(��y;����+<���V�ܮ����z���Evu:��2����=���!�K�[�xWK
�il�����qn��>I���-��UI�rub�j�=Qut9�{̝�#� Y���r��q}�V����� q�n��6f������O������e�� �b����`���g��8t��A�ש�x)n%�W�7'��C]$�3�������M�s���-|��f��9��A4K�l��@F���D�����,��ߜA��[/"*����%�="5=�He;�^	1#F�,"�e���Zo�^?TV����_��z�^ЦE>@�
>�$�RtF��1~vu>'��s��K��Wk�pϚq���A?\7�~ϟ�_�G!
����&h4�[���

d�.����g+�񿩧z�N �C+�ޛoxt��mS�j�����;�'���kpڜ�L�]��)V3�� ���R"�@(����l��t�O�;���;�
Yͣ>*'�a^9&۫]�g�7p�v��W�&�C����C�ޮ�����lloP�H�l���(�����X����}�`���cZ��S���h݋�e�9Am3�P�<(�L��ho�|�h.Ϲ�о'C���F�"�ʉ苃��7�Jpk�xsJ�3I�U�X��V�D���6 �OfQ)R�R������r�l�i��Q�u�)��-�a�5���D{j�b���5{f����컈@����㠸.;����}l���p~�;(�:�6���,�y��{?%�9민
�8=*��I�)is��c{�{�#diۥ��,��lhq���W�!��a s��[q������%�U�?J(e(�T�sZ�%�����>��RnӺ��j�ܿPs�>��l��n�wEl1�u��O�!D�	B��Z���bC�~�3Px0{�#�PR�_�L^��,����A�ǁG�	�?S�א+}�PK   �rZ���7z  �  /   images/be8de2bb-09ef-440a-a2d8-19619bf9d0dd.pnge�uP����iv	Y:X%D$���e���T�[@���f)Ii�R)ARZ:�����>����s�g�{��3��+Z]U���PA���֨=�A��U83�t�7�@C���o�����B=������r����p�A����|���ae�j���n�u(J��FK� ����>�&j� ��"�>ݽ���vЦ;������p%̑���a�Է���Z��R�P�Źy����S�3�g��'iĞ�j�8�Z�%�Ww�G~ڝ�ջ��\1��pY�ӭ�Ǜ����L�>�����֣�I�'99y���������_�_�"�m�g[#�w�G��,���o\��%�*��&����o�i�7L/�f��;��`�Ҳ���>r�92��{�H$�s�٣���<??����QИ���?��)�G��5���>����7��II8 �_��ia���0-��;���>������r9�ﵗ� v��eE�|R���k?�-?=�l�o<�Cj�A��Ӳ	~�e�t��w�´������K(�
�\���.?a�D	�:����'@7ݬ���� ߽�����}aG��o�d5�J0�#�I�� GD��i��p!�X�x�l��G��@j>lF{�����O���`�'1�		��`kQ��k�n�+�߲֕VR���@H&����ѩ�_Ĵ��� w����[Tx���F�s*�m�E����N�*�]cX|�<���"�P\��҂G����ؕO�i
�=I�Ҩ�8��#J�h�6:N/-��ڇ�-N� 	o��Y� �����O�E��{�
�/���L�kp@�wy	d�Dލ�V�����M�O�ru�Ñ���7�M*�P&�i�$g�P����ơMؒ�?J�x�]�'6J-M��%	т���bq��6K*e'竏*��ӰM�%����[��w2��S��፮E�@y7�J`:��;��Є�>�L�Jq��1x��J�
�O��[y�mN�P���].�H�ԋ���k7�ܢF�G�u��`�e�Q����<$��v��a]A>4�6t��J�`���&���7k���sJ�=%Nm��	�烥��+g����\e�tC}ە�nsߗ�բxy9�WW+�IfQ����ȳ�ID����)t-�=	�(Ke�z��+O/L8��0LDQ6�P6�(�T8��C`�)��ڔ|Ox���˧!Y��u��`���8���[�}��f�/�\��S���8�\�����^���B���İ���B7[�2k�L�t/Ũg_1��ǃ����p�ҌI[�A\����&I��ϸ�G�������4�ihI�	CX8`�<!�����3���xnՎ}m�}��Hui�!�6��ޟ�^��D)��_�]��� ɴJ�+Ţ�ۅiiC��
_�$���b���BF�GHā3�%���㘂>�{:���,?�f=�i���$Ga��m�Lx B��Ha���8���݇�ǣ�4_�(U�&���fY-2F�'"�A�^Ui鱋�lB�!具�"ZX)��חI���r�6�9y�@�nj��Y�L��KvQ���� 0c�'�[����ǘ��1�ߔXb� �ٙ'�x�˓�q�
�b�������Hά0�A�8�.���nc,��|qrZ�ޖ�����+Gٽ$]�6&]��L�u/,d7P�����O��4��rtQ(�U7���[PX���Қ����t�����cp3�
͵\Q���l�;�n"�;����p��y��!�;����Zt�f��>jg��ƾ=��O/�^���TY�� `#o���t�L���QD�����-��}��B�M��es���wh�Ϻʩh3im_�6Yb���lc�y����]�0�Cw���0"�M�2n;��85{���Mݱ7��uҵ`|%A�z!}���
i�VT"�X��e>'�}�	ռӲ�H±���l���b}�?W��qɄ�������E�W�M |��L"�!�2WW������tcPh���wDpo�F�P6nh�����[���a}��I#{^��X�p��ŌN[��j��*Q�==�%<2���;,r��$���7��_�k��ƚР��
ݪ�Fs�S�}[�|W�eG��������~�n�"Do6�K��u%����a�E8��F�D|��2��C���5�^��q������<O���ƹA��s��(��4��(gp���9U�0���޳���TTFHQZj���z�`�k����	Y^�-e%�ˠ���܀Û�����Dq{y#�r��G9�2I��"�Ke@;WҪB�y���hF�z��TL7�&�ȨD5�2K�> �Z
8�OfQyw�'�!�2�q��-o=lq�E�O+�˭�X��'n{�^YOI���v����y_�V��o��)�\q3?Kf���^��T��l��]�Tӯ5�Z˗~q4��#���W�`�����Z�������ed8>%�Y)-�	� ���'�;���$g���)0�Fǔ;`K���l (���y���S��O��߼�>��r�sQ��l6<njڛt�!
��<[mg���s Bude��g����1�\��"�}�&��2?���'K'"��/$b��o�2v��j��{���y�0j��C��3ngZ�;�6�`�ݜ$;��TJ1>�jll���8�6a,|��F�]�ٹ���۟�;��V�Vqנ/���õynG�jo�M�+�ݧ§��~��'��I�4�^O�����H��/Qδ�!����jz3�����͙�b=6$���nE�{��k'v��s���)���`�E���i�g2#�C�=Jj�MO2�����z�֡�?h��F��8��y�&l~�R\-h3U/�q�������������K�h��|�����X�I��r2F�54H'��O#(�Tf��*?�و�����}��"%�����ۯr]�C{����T3����0��6��{�Z�h=��~cdr�go��Įj����g���3���f�z�g�[&�GՉQ[. �WNn�wU�o.�#P����$t���!� {z�ѐ��s��L&�_pgk��d3��[��]p��d�*q'����wUN#(U������~o�0�����g���J8�rC�@g��%֤K}a�( �؍�Vy��%V���(d�ru޻�����q;��]�J�W�a�~�&��L3r�a׫n(*��l"9����t'0�@�fE������t>���Uen7���i�3-�7Hw�Ol��;�����L&L*�qLoFJ��?dǰ����H[5^(����+1$=�\���e�9�L�^�^b.s"vY2�j�|�Z��6y�n�J�E��j�i"�����kd�|��"�a� ���J�����B�F���4d뢦@;�7T�K���a��x�Ǆl��!y
6���	�,QjK�f�3�	~�X�)X����K�[�h掲�4O Ϸ���V]KV2���<�/�pn� ^N���. )��r�׀AᏉ�<�C\Á�}���Z���G��ˀ޺����v�N�"�W�ȅ�؊���ʎp�&{������*p��BZ�!(���������(�[�S�13�i��"P�%$w�Dd2c��[�k�Dώ�ǚ���ux������`�����͇����Q��
�4�T�f�k-���;��)����^��Mc�*���ggҊ�գ�n� SE6N��n~�iP�/�[q���ʮ-v܅y�R�ˮ���뷖�����efx��C�N���ɽM�O�gq.?���ֱ`�ь�ăz��'bSrԍ����to�7#���F�a/�C`�e��V����^ZF
]~p���6q��$r�`��$`�@��N���y��%5���#�P����ڬ^�C�q� 0��)S��2p5=�����d2���g�Wb�>C�&���]�Fހ~�Hl�G�����!~�UU�F4��魕��]��#�rNWN��r�~E�Ԁ���x����ݛ�:SUB�+�*Al:��}���P\����1���C�uRO\�K��X�}����6�be�~�ܶ�_�x��8y�iL�L�\�^�܎B1s�,<o'��=��$<����(�a�8[�B�Qe��c�3��4Y�Ҧ/�u��	T<?�N��F���r��|~��6X5A�H�;��5mЄ�Y�޴�m�A�eU�9���VtU���G��{ؼmX��6���tT��J�m����e�x�4�Mۇ},�n2�H�.E�����ʥ��Ftv?���f�[��H��.Z�;9j�Z�����t��~����e��V�K�*ߎAq�D��,�1TP�Fm��c�
��z-��]����6�eX�������l{�U�=N�u\:�M���]M]�T6�c���(��:<&���!�w<�q�� �F�s
�6� �`��|ѐ�
�����L�����qbЏ��1w��;�i ��7:Ќ�_�?����B�{���F-�`d1AcQ�o,�b��Y 5�d�{��A�l�������;��_�U		'��=;f��?�U�	��5�|��������oWtp�F����t' Yi���g��4�L\C�[�r$�	n��4�F��μ4�;h��ޫS��W[4�[��u�jX�>uW����G��ٯ&���ۚҗ�X9�?�Ur�<�6�O��'�[�F��_^Vj�)7c�1�z�s��0�����oRrNq��t���f�8_Q��2H��q$?��AY�j9��p�_�{�U�6����-��DMn�u�z&?�ϸӮ�dk`��Ķ9��_Ā��iA�5��yv����ꋶ���M娖~,.��^�gį?����J�a���%Yz��v��#K˸�������*C���}�Hx�ټr:/����\��,^�A�y��n��k����>^7�t�L��'�
D':�ϒ����/oٺN7�]����}�j,)Ѿ�R��ɲ�<�2"���	Ym=�pXG��-IgN����KT�lukL�>����L=�Z�zAC�D�F��VZ�q*��'��������Zd���6��7��g�M:�7^X��Z���h�!��Ŭ메"X������x�9A�6�	��O��4
e3���h��zDxg?)��Y_�(D���,49�jN$��˚ůE�C�	g�Qe��f�{z�0j�Nr�̡�9�s?j@Ǳ��Ml�����C\�n��{��9�ۡBھ� 
��t}����|��Bl�t$�#7��57���~����Q� Ll�d��ͽ8#� �1S�_?�1p���������-�JZ���]N1�Wߗ��9�pP���@�?Z����3�U������H]�'��(5�F�kx�<�@���qbM�qZ���(�����|������i�A�n�<&D�V��̒���x%0��=���u���y���h�����kӶ���K��v����yMc�t��8ZvR���֪z�~ń'��rb^����w��{�$� }�i�R��*|eciN��<`��Z-����0�U_��e�3���K�s�֠W�]�M�%�hh��)����fO�3M1��b)��?�]��l''�M����sTBKӨ�4�׵�j��
�����9y��ऻ�����j~�iF�T�M���k��>�����3Wo�`A:�FH����X��p�>��
�/�ii̮����g�DU<�&&͚��L������,(=��+F�:�E�,�0]޾8֗+�_<b�|}���u����X�^j���cL��5�Qb������Yytl��k�ǨLM=��?�/wĉIX=#t��qxG"t#��*ΟY�]�t��7�1��_#җl�U�S��q����d��g&t�znn\��{,!�)B��q�P�P��p��K��M�	��޶��C��μ{B�ZHR���x�X�OS^T������9�x�sS��$����R��ǹB̬��F�1>z|65l����M��h7,��>�ٱ��2�۴QBb�(9Rz����ϲ��>���e�������%�z�8(s�IS&�/hDu5��o��r�%(Z�
���;�ρ@�S]��,R������ڬJ��@!�_��4ƒch���%ѓ^R�6ihJV��٨��{��`��t�\FΥ�E_��+�le��_�o�E'��V�MmE���B��������5FClwh���&�3�;J�K��X���HM|ląv��K��D4y��-��������[�V�~���<Ź�@����7�:I�j����H*N�W%J9�P��O}Q�Kj?�Ո6l���>݉�g�����r	^�S;�~;"���Տ��z�n�f�2�����XBDF�ڦ&Fީ�����>{��58�QkH�';�:�1-Clx��t��i��)W�X
( i�ޙ��2�Ow��9?�׏��0�-G6bdN(�����7�Y�~�{l�vz�������mg5\�#{�����0�N���3������\F��7�H��rTD3S�~s2������:`�8�ER�,�;��[���mtܻ�ݫY�!��w2CS�ܻ!�>vK`���Uf,�&��xH��,9]��c�b�h��R{���8o��K��z���
�y+I�Z.t�Ӽ��:q~W�Pzh�Ֆa�Bɻ���
����+k�]�|Ȫ��H�U���5{O��ǔ|�I�͡��^	��Y+N2W���"�S���V-$�{)O~�����g�;5��d/"@���J��W��txnh�EU���Z��.YL��<G�3�
'��!::�'�J��؉/�Z��F��-1�͸��>�������M0BV��ہ#ׂו!����|���D�Ko�<�EY�4J��mZ�5ԓ�n*��R_�|LMܫ�\�Xr���(�bx� �(��SK��t�2�|�x��]5�Ey�KI�i��c�A���K������������=�	����h�U͡����*�f��� PK   �rZ6e�b�  �  /   images/c0cd0a79-4e96-4647-8bb3-400a2b193618.png�YePЦ=�8����<Z���n$D���H�n��n��n	ii%�������ogvwf��g��_;��j
�x4xhhh��Y���wp�Ÿx|�	�a����������h�+R���k;Y�{��Z�yyy��stp�0s�z��j�y"A��F�(+����7�R���4�����j�����0���Ā���K���%h+˻���#�����SH�L"��8:c��X�d��˦��~����F'O�絍׌��~W��z�7|��;����d�CD(�Gg����Ȅ����S`s[ �OME��%��!�HK�VP�'�M����<���fU�*6��(�1��LH����u>'��?A��3, K/56���'���W�er`	�<5�WåvR���,�Du�b%�\Β�Q"G�Ni�p~ⷄ/��0Z�a���3Q%�`>x9�e�1#�b-�X��,�Mp� /�ɝ��� K�C/�*����&�U���oґ�9�N�#\������;ɼw֠u�PO.�s�V�q�K��= O�}�)(IH(q77��En�3���&���Z����[��n�:�9��İ������XYܞإ.#S��(CR2��Z�V�BXp�Ll�#M]���a�
�-f�*�&�үN+6h2l��Vb��9�"�%��Iʿ8�}NFA��友_p�V$�n�-B=���į+�����"��>aH5ğ����i����V�:ܞMpi�/�%�������0�Bh�I�e�uv�8��y��.*M����p��v�Bf@ 4�۶��u�uR0�f�JQ� ��Ǵ����\fZ^�9���7���#ps�:�֮F��*�+���g�M��}��D,H�����Y������W��;����y���#4j�}����>���˶�Z��g�K��h���Rǝ�}��dp~	�Z���=�)f�9��F-�g>iCb�4&!������&�ֽ2�����v�
��&)��l���&�(�	����ƯVjzo��2���{�����)Q�z����e�GU�����nS�US����6y�j�h������#k�EY�AE:r#��N������&h�U���q-�^⑼���ԛ����ԅ��I����~(���Q�T� e��0��Y�5�V�1�B�F�mo..ݍ����#;���>*��Td�rb�}鯻|��~J�擕�,��\U�P"^N������wT߶
�����R@�����9�b��u�pޓj+�|}�=����W/d��n��2os.�E
�k=+Z��#dK��)��m�L��<�a��gI���*^�"��R<��':�`���U����/B���տxNsW���U�N>�x˒�7��I8T�\#��5Q��p�g�4�~β|}������+�n� L��΅�?^CV��r�q*���6�Ⱥ_r��4��ѫ]�jIV�9������B}�((�������w;Z�ƋJF8��M�S[�Z�b��������,����Ju��=�a��,���ŬD���^-[�9�[�u��]�ҏ⫃�"���G��er1��&e��.,xí9�z
q��h�ɰ�i<�G ��0����t�/w"m?`M�,�m+����T*J�]N��_��fw�^{u��|o>vO#���j��Lg8���d2�&�Z��b�؍0V���f4 �~�h/ͤ��
_�{� ��A�I�9y�����B�K��L���<b��o����^ZEC���`�a���?X�5צ����b��K>�3&�.�
k��C�K�=��Pּ̑��j��a�RqF.�ZFЖ�-�ΦnZ��v��*zy�ag/b���@z(����l(����L�R�E�8�7Ȗ��f�0�9�nk\����5=^�����>uG_���?y<nP�@5�9����jw��>���a�6�Z$�?2�ß0��u�qB����;��x�$�8��.�sFy#��Z�C�z��R�
��m�#B�C���/�p�!� �p��c��kbdl^Ϭ�'�h�u����@w��G��q,�r���5��6,5R�w��������!A���Irܯc��A�_��y��n���1+�2��"�C��Pb݀#m���`�|�Hf�����F M�c�7vQ���ݏ�I/"C��Qc�3v:�J��:���j����B G?L{�hP�S�9,�oc
����w�B��/3�������J�ˉ���l&W\`�={�'
���]Mc���H�Z���p�OI�F�ۇ�[2�)��u
���&D��x#l����Gq�!*)/�*�qK�I��*lq��^��{数s*G�MRϿ�?4���(���@rs�s��]l���f�Xy��c�R�F�������SiC�f#�?2ښiZ [�,�9+�$jw��i������LV�	ܜ��'E�
�v�!"��o��}*<�Z>Z���0�l���2#	O�E�}H��d��
ta}�����	�����p��j8�����έ�8�4��'"��Ӷ#'�zT�!xY�6N�,n�1^PL��]���}��\�����1��)����m[�T��N[3 f'�2��[��:��S!���`%ۢ����"���"b؄�����"��=�N�BC��@�%A5C�:�����n�Z{�qM���?�2�Q/:j,|�w�f�6�.�-�f����l���:Sh���E���K�fg%�A��y�^ǔN�e�������U�k~��0�9�1�x�\pѤ�y/�Q�\2M�yrn��X�!�xG$=��hm/�`^V���Оq�w}��#Ǘ�M
Q�.���u�+]>��GQW"����SӐ/�!)b�|�n�ʹ���^�T�D�@��s�D;�sN��L ��s������hHA����r�N�u"VN ��9$����O�����x=l�f�X�I�8fWē�[�|�����Q��V�bl��%�`��������Y�&��4aon�*�՟|F�Q}�~L�o+���_R�#��'Ҹ&��-�#���L���'�����fW��ķ�!G�4bK�8Y-D~z]�v ����Y�ˆ�;�=^�װ�����<��n{�)n����BI�)���ltm�{���&'&|kӛ|�~1��3g<�
Aʈ%afs����$$xHl7��|:R������FY�6Qu��)���ӡ죢l>:��*4��?�bXcF�86ԏq_Q��J�KZݍs_Yg�_\��N�.����\�;�����-)���Wn��M��lgӠDjVT.�痏RěA��mk=�������T��>��oE�U'�6�ȖCLn�Jy�辶� ���� 	ө��a�[�[��?.�=�s�mp#��~�n��io���٣���m8�9Ɇ�GMD���79
&�ۢ���,0!Gl�ݝ^3ɕ'h�����]�����'x�
,�Uܕ7ě�w�wr�!�ڌ����z{q�\^X��Y�E��ދ;��[�p!m�����}�9��ˈ�6D�7��E��_����A��.M�p~�ap�~$�S̲���2W�}�7�X<6v5k��w6g�&����/��H��leIHzj)�Lt�fr�ۙ�ͭ#�+�o��������kԏ_����k��S���I�� �lVл~�>��Ͼ�]��疽�/��m�x��7=������>�-�dB8F��*�]� G������șUIT�1c��'>���������f4�fq9	��s�ҿ��d݂�)���]y�ELf:���(���tP�����gn8�}}S_u�JϘr��|�=\�P���r�oRE�Mo�pmm��<f��L��'�g;� _QSc�v���TFbX��G���ݾ���3[��w
���V�����j}"5�d��`9�x�&���Ϫ҂�j�i�S��_S� �g��b#.����!����Dy�9�rnyԶOZ�����;K,gR�2�T7�,���o���RHQd;���%��l`��z���vZ�ɴ�J>��#J�*�v)s5�[��o7P��
uޮƺ�f�pk	��{��;�Q�TR���(@������ę�w<���њO�o0-ȁp��÷���$��Φ��0�J(���ګ��z��/9�nD�_�j`:� �b�j��3h>y�5E�D��2Me7�.��np��ޱK���I�u��{[5)����J��}��O��-b������&C�I	���%�)��jן�\o4�1<Rj= ������z����K�L���uH믒�"�^�g� S.�T� 1|V����!LPv�!��$[ 	�������Tsy��WKvJ<�aXv#�I�t�H���`F�[Qz��E�n��`�L���m��PN�AAQ>�"���`Ѳ���36��ˏ>���f��d}j@�D'{�/h<�c}��s>�q�/�6�Q�:_�����df_���������P�&�:4��g#�����zx�(�>ҥ�X�w|����|(�"���*���R�g̛�>J�B�Ok�oD!�mH,�/fW:X�^g/!���]w��-wT���Jn�}Ja��2�~�f<����:����,�F�w����c�-�Ѩ;���*���s�ڴWf�zC�!�oQ~9��(����Wc�>�9Ue��T�%l
���M� +�R/��f���#��|oÈ����@��w:%FEi9�=�u���c�ceh�����g�9�������F5�p ��5ony��Ċ�ƑX� �I?��Y��<�M��O����˺OO|���N�9a�-�q�0��Q�ͦ�+[�k���1�����i������=۪m��M{)͵�uV�7Ƌd
�*8�hF%p�!�Y����V���Y9�)�����7���]��ޛ�ݮ0�"�0�΅p�z�R��l��+�Y�>����3W�D�����Q#�Z��e��i�05�Ԛ�ì9�� �R��������{1iR�8�wy�'�'��8�
�DX���A4_M�;�S�h��QY��}�e�#��-�m�X�!�V۶
��1�M���*Hj;�D������KB�O��S8i?%߼��MRZ��m�E�q�`ʣ\m�K�#>?v�[�Ռg-E�{f|%w9�8Fu�ű�����K�� ���c�����J�xhM]�e�:F��G�1HL>o���c6���e���a�{��aKL���鹲�Ap��8eo�� �������]-���Td 8o�{��M���q�c������-�p Xp�Lp���~&��ʭ�Q:psk�����c�Ui�/c��$KQ`�x�B���ϟ��?�:�8���܍��>����<��� ��$�Ga��D��O+������WSD�,��lCNP���6�7�ȏv���L��P����gxE&%���������S0zS�)k�%em3�
���M3�z��[�ī3�r���{l��1���hp��ՙ��d:���j7����9-�C�"�Χd���eߣ�z�If&0�\�/>c�BW��|P�x�Y�[(ɕ��H^�?���	�M'�������7?%ݽ�j�3-iW7}wX�z�.KP��{@�t�[�QC��I����,d�<r��i�7^Hkɹ�>0ا��ȫs_&*�~�ZQ���־�����=>�z����*w "r/`�=_��?�}��l]�R{i�x;Q����4J�Z���3\�����jh(!����K���x��
I������\޼� 0��+���	t�$�#?BzF`��3p݀��o2TT���$pKt�&�a�
g]�-W$.�����Yv��G�����������0������|d�qS�E4╬�3⓱6�ڒ�=���:j0~�l�O-m�C����ҺQ��*VZ��n�'�FQ{���\ld�B�ȱ��Q�:��+KT~�*����?�w��lN�:�c�Dh��Y����y�J����,$���Ǔ}`�~�������C;찤Ƕ�#�l#��&
�{����k���%��N"���}cf�df.�,�K��#�>�g`Fv4�O��9��x�9����?�6�?0o=;R��L@�����������?=�Q�a�k���fF����3GТ�r_�������@��:�u'��"��+?ʳb��x�'������#����C�a����e������}p����$���͍��&N���v���s�;H����$(��贒!�������FŬ����`V	l�K�5V��� 4X�G.~'�:��H,�9�&{�5��L$U��m���3M���빮�;��I��y���I���[}��1���;@���#Z�
���b�@�8��J{��=.�Ѣb�.G�+���_HiIܸ9�fqe�O�ߣr'qx�0)�p5�ʒD���¹�Ⰹë�Oqp��c�U3��Re�F..���ߐ��k��/�0	V�Jּ�l��~i<\��̼E�paTT`�L���W�
 ߞ��YK�_K�Ǣq�S���SI��a�\�,t"������e�ƪ�jGTNG`����˫�7B�Γgh��\'F&�^�/�D��˽��%5+�GE�B5tM�'���a�GXh'��s����՚(pFZ�I����e��0m�������?7���M�⛿���;#cU���[E�z���D9#t�1>��;�o[]�=�Rн�G��02�3P�`Dh�v��f=�Nl�:�^g2�������:�:������S`���g*w>I�%_����3`��RO���*�cl~���ơ��}إ��閍N�eg{J��N��Q_3~3�[��`���8���@i�";��h�q�Oov�:�_i���m͉C�k%�w��ǹ�&J���]W��k��b|��#� ���ny�� H��];.�
	��;|�}�eڽ��vV$�&������H��UĮ��c��8ꡌ�ߥ��GZ|� �*ז�N�)*�j�"'�DI��!t��/��Ƽl1�#��j�(��ي�ǧ��iY0]|I��C�#���}������;?b�(���r��̊��~(M����G����W�Ȉ��N�2�?��e:u���9H���E�u�ƲGO�_�1NV]��^$P	�7�[y J�Fb�(Z��Gh���� �d�W���-��A�Z�Їe��G�>��Vϰ����C��h�^��1q�%փq�5񣅨�����a A�9�jl��tflR���b����+9I�3� 	�$_�b�2ػ����M��Ӊ����wK�i<��7�~��yɜKR�G�1| 6�P��ҪotF��TPS��P�ӌ��C	!��i����D�X��y��>��M��ߋ�h�U"�,z���򭁏&�=U������.�2���AW�Ԗ�g�՘����<5w��i�\��H���6����?�?S�S������PK   �rZ;mLF   P   /   images/c560fc9b-7045-4fe6-9a6e-de67d6663603.png�yuP������ �KI,�tw���t+��K�����  ��t�ҋ�% ,�-��S:~|�x��̹�̝3sΙ��<�̉��zNBDG  H�e��~�00���z���]�������7�x�uWy��r��xo������fe�b����6s_� `Z@*+x��"y���'e�vT�a�B�ɥk�iB����/P����<��G����Z)������5*��(X�Ԍ�������-7����Ԇ�a���_�ᭀ��)m���8cE��Bdq�S�� {�ޫy�9��	}mQu � �&0��� ���B��z 셷c�	�¡R\D�.A�X��K�#�w�-�w�=�}�F�n�M8�W���,Sr�~\�Y����{/}�y��|j�Kx���� �(d�z��^����Sl���;UH�Z/ʑ�~o���ˤ�����P�R���V�Q����W��9�L�z���H^�%U�O�],x-���H��+����-w�m|6p���	�m��=|�Zhn4v(+�ȑ�ǎ�����oOߜ�/�i�]�|�^��o�k��<��6�R��؞����c��v����4N�n�kL� �b��9�w� �������</G������-5�?�[xZ�W'��?O�����e�?�O�!Z������:m�h��`3�8O�5sU).)}���'m��� �t�5��ڦ�1�;{���k�N͓�8��쉌w�k�Z���Dߩz�9qS-(��__��<�d�һxwn)��\Fr�wj�����w�[b�&5eN���ӡ��4��C���N��ƍ��v1������$/h`��$��n�3�?������q?��踝�����MM��{�B��"^^V`��)��)}��X�ow��h"��	��%8��7��Y�ʟv��6e�^	_�+���'p���h1ʤ�zo�)s3�n���2Lh3?��������z�$'�LH�=J)�
�Eg�宱��t��6~�EeyL	V|k*������:x{��d�A'+�H��
x?�d�Aч{����El?9��>��\b�cs���wg��
؇��)��k�q��o�ϓ���Q�(n�q�H: f����2�L:=�w���;�'M&�92v	Z�O�g�CH�h�Z��|���9�u7��c^M�� �k���eK	-Z�����%���`����+-�R�p��Wx4x��=k}u#158P`�a5�!�
Y����?-�>e�'���wnY�n.w3H�J[�����d�{��@�jh<�6�Y� ��B*���o>�j�C���r\�pt�ﾤ��E?���*z���U��C��@n2�`�b~��)��-���q�j�)�
BpQqO$�.I7����.��^/��]X��W�4|ğ�d^ƗI�p���'�=����`�n��{����r��9M �>�;��"�V���|αʉ1��B�4�M}����������td���:�8�3CX�{M���f�[�%͈� ��j��y�;XUxu�m�ЗT�1� �U�'�EB�:��6KoGFӸ�Fw�^=�3��B4N	����=��搉 �v��Uw�j5�-ψ����@���x�qZe�������p�6��V�>��rF�QQ�֤�j�ֽm��%6e��\U��4�wb��
Bٽ�)�b{���w��rp#Ͻmj#�� �qMq��M��Nno������G�\�to��h�?N��iʧI�,���(��/�BP��|��抡���n��g�u�F�~DYi�0ew6[]j'�Z��G�
R˻�K-a�BP�G�.�$1��o�ď��4lBi��Z�9�����Uq~������&꩗�oB�Ъ_��`���N��rdt�4��F�Q#����@,3��*u��]�c����9i���}���8���v�&�t�V����d�%����Շ0m��6h�u�f�ȕ��Z�zQI�b���5�u�W����Fm�ԝ���)��!�4��L��K"=	�A���o�n a�Y�>z�*���C��Zuu�e�y9"co��֯� {��$��[�Z�G�D�"�b۾5�7�Z�M��m?���pdQ����n��٠��=����_޺�a�1>�����xl�W������̿s��XF�_=�cd�Ӓ�E���mϿ�keX�U�^ ��fQ�N
�4��J�����!#mz6K��\X뤵�͇ƛ�xY V �_m�F����0yID�SA/0Mk-�v�
�qu�Oh/d�='��GÎL��0����ٻX��
=�PP��o�w�<���@��=�;
dj��ϑ�=	k�O�/�zd��=DG�iZ���J��0�Anrf����:���ˏ��W�<�ld6�v&?b��_0kz�۽�y�K&����-��R�r���#�c^]ӟz����e��!�N6Xr��<�
=��K �S���p�vꤹt�|�L� -�S^xBS�~�0�b���8���1�q ��p84L��x�����ʞ�Y���aY&��r���;���/N�v������hW�XєT���ǖ���x	���*s��^@��G(T�	Jt�<p:�M��;��4���6�������
�1H<K��؟���t���CO���$�1v�l�e֔@�EzLu�8@c���=� t9W��E�$/����+*�:���9�}��x釀x�3cV$��R��׷f2�D���yS�y�xrh�~>fp(�C���$�� �z\Բt�^u���`JZ΄{���Z?3QR_SC�b
f�>���|=a �$dG�av/q���wvc����ޣ2w��at7�Ž'^������i�s��$�+��E�X�"$;m�5\�4(w&ѻ�X[�p͖63��n�x� K�ހ�ڊ�դD�-=�:�g��~��G�yEh��; ���U{����a��O�|�����Me��m�,qmD����vF�YZ���HG[�\�7'���R��1�t�/���hړ���!\2�9����4��q�L����Շ9p�A�{Tg}�g�;U:��a�lM#3FC+\lQlN'�^�7���z���\���n:v�B(�n�������56-�b��e8_c��
�<���[�}��B�[Z�~DHj���M���#O�[����L 
�H��#�dD��Ɖ��6k�y��<��|�2&2~d�34�Z�x�ΐ�krH�L��� �ӏh��}#� �ui4�W��Շ ��`z]7k_�e�E�g�*"�\[�E�Фw���4�2P�2�Md߅ģ���P�'R��K�m>۸�U��RW�4���i��d�eN4�d�o*aĜ��{���PQC�Gv�����%c�Z���Wέ��eo�ͥ�b��r��im����M�)�������X
~T�E�y��Q���ʦ�|Vѭ��Z����P���^�ѿ)�������5C���lЯӋո�?�g�PS�5�Ɏ����p��T����CQ�,�t����@�8��OC���&y��!2I���(n�hV]j���yW�Ҽ���[�5�E�=�l�q���ڛO� J�
r��V�{L�yGl`k=ݷ8�c��f���[��.�� xu���J�A.�)c[ɤ�RUc�\�t|���vw��t�K�\����S��8�O�=��0Nh�y���(��Z
�۳u�@)���6U�Y��W�����Dmܜ{�2�֣Py��3���	q�4�E��Ƽ��5ɷ�U����0�@��7�`�c�"�f�烥�������=�~�NF�9���_mC�s+���Ƶ(��B�h����;^0������q�BB�5:�D�I��$m�gG�������3���m�?�x�X΋`T��]r��a�3�O�ͺq�]����<�"'i@0%P'�����c5D2?��u�~_�ZjRȹ���J�-��)DbY���.ģ��k�۴+??��U�����;=�_/D����A� �{D�b�s	j�Z�Re��:���"�j;?����IM�ƥ�|v~q��+B1���s��mZ�~D���[�Z�6'��=d���_1.'S;�'5tā!qF�|�N~�\�Yr�Td��޴n��3�/�b�g�CA2��c�ԅ�s!V�ƅ5[X2��9|��W�������<�n�v��H>��x��Z���F㶫���o(�
w6d&�F#)�2"���Le�$0�R0�	-�DEȩ_����5��U��`!�]1.$����^9�0f����5hs��9aW��8/�2(���|\c��ꔛ.ũ%4� �mj�����j~_���� ��1��]�?q)r�[�sS����[�@���;w�|��b����],��M��I���j\���q[]�0s��^| �X�U���zD8��rAN����N�|�
�˥�����q
��]�ת�����%ݩ�-ł��
��4���3_?�9�����+�`���I�Q^�SߖhfnL��k2�cϙ��4� %8r�{�l-��U{'U�_?oc h��h���������8�����k�m+��A��X���o�|��z:s�&hIǷ�ۣ�ůȤF�|���?���<c�$mq!���轭��:��kx�~����0ۧ|i�oV٦q���������c��?| }a���/�`16G#���xW�65{���-��iU�H��U~ɘq"�X��Ή��G`�OG��
��г��$��
B�҉B�9��iGoR,GHb��S�j�Z����d'5�gtI�e�6�K���8|�H7_0�m`��)��bg����n<�{�ƭb^��+@��'�����3o؈4��|�:�q���3��i�1巡�u�\ɿXk�id}�>����-�CS��g���nl̟��|����N}��Ko*�e���։ׄ�������ĉ-��4���P�E�a˟E&x���|�M
1|V�^�n7�@�0���B�ߵ��8��l�m&!�4Ӡr�=+_�nš"���m��D�ڨ��c������SU��#x%�I�*L,�/�o_zUSj�M��6�����x�\	�cOI��fg�9*6��.���R���� ��^z�u�|Kn��M��2���3����r��u��~g�ŧ;�{(Y��9��_�� �p��r䖠#��� �W=l��<�}����%!�,�	"5���5� �J��$׶gC!��=DR�C�(vv��@���(4Z�'	�o�TJ�~o�ٳ2���`a]��1�y(����U��%2r�eɋ"�碿�8OWt-�]�RƌQE_!͠����F�i��g�Y�I��%Ar�o����`zi�d��|O�ʨ�}0�[[���8�A5��!b����oUԭ�p�跙�/�5�g��skf�Pڤ�疔͍x�����ѹ�ʯ��F�o��e]g�+���KDs��c���n�W ��G�{����S���)�_?M&#����.��s ЈA�B����7,�z��gx>v�� ����c<���g�N]��@	9|���� ����?�
0�h@zi��ho 5�b�O��34f��*�13��	�
;�@�<�y���'6Q��a7.q���m�]f"ܪ�+D���uB��BM�|�(0S0�3*��PK�`�QZO�W�ߕ)�'��>Zǫ'�&�NTQF@�4��ଔ���znW[%^�u4|Fcpl->��X��q�r�����3lP�'��(�p-��� ���yb�#&�:T4�&'���Q�xa���GO�BS�]~�]��aӜʭ�_X�AĆ��s�YS��ɏ"������
4p����R�ܥK�X�nb���A{�����)�|��=�%U����Xr�K~��i��`��rʟe)�őSi�AD�)c���+�w]�e�Q��w��3�n��Y[�Ρ����>���):���Ƣ��rX,��F��&N��O�m�Y<�kEyL�,�2sDRqh�
8�G"�^�a��	+�6�W_�.I8v@�
>%�9��G�:��C����O5�"���/��8(	���j���WG��ۤ��p��,cjKG�l���M`]�6Y��ʯ��̥��?K ��rA����%"�������\@:�P�H���,���7rw>���-�E������َD�U�rkҺU��Ex����ڐ������Z�^=A!�$��,������5(NBl��=rܥ
Bi����耂��r\�{{$�Tـ֘�Ц�O����:�YT,/��ד����ַ]}µ�5���Ȓ� ]S�>/�͡���"ahE@�:ך�^�"�F�'�m�Q<CF�(�m]|C��t�?���#����k����j�K��C�^���@^��p�s���u%�J����P[A/-:��u��|�ʱ�V�Q��6Q�2�@�tY��-%�����sԫ�!m�1'�늇�`N�Z̮�f��D������۠��7y|���+�쒂b Sj>���&��&J��'2]���ɺ���AaB8��N{��R �����W����hKa7�B�`�@�)�=�_��³�x����_B\/���.גH���=����2&�U�7[Ԋ\�y��:+e�����'�q�[�<�_���ln@��X~,C������`6���%%[�����*nP	=UV$�[���)�+����������`��f�q�!)0랷�ۢ5R�b�LyZ���4��L�1���ĥuj��V:���J�GZ���e��L��+
����k�z��ҹ�N!�]n���\�@�'*�ߡ�I�a���8�1S?Z��>�s��^���\��0�4"6נ�g+��;�z�7���X�b���䩯����� `'�a�ZDCm�{s���Ҹ��L�p�nd���	4;�a�xi<c�ة�K?�o\�/��ȁmG0��< �?��n�ݨ�G��ݬ��@��]^�w#�B&�� ��`�|*akI�"���8��V@�V��IS\��Эc�CT.�z]���������\q`���\����Hh'�Ժ!�㨛���8����� ��O�С�����5i���s����RuX�%��V& n�����K����I(�o�!e�N��=�y-J�̝���\.��M}V�HY��Qf�BB�i���2k!Rr��W����R��j�:bdp�0�i��TS=�Y+/��~��KȰp�2�����C�[�u ���*�ő[��f�.m�G�	^��Wd|��d�g_@��|���g�	�b�+-v���ͬ˭�t#Fƀ��]�x� 7o�˞��	ҿH��s�jz�ϔX0����,�0}���v8���2M���i����ig��[����G�,'�"B��_)*�4�ܵ�`��D��|7=�t���~X��0^��S5~e}��*</&�̶By��y["�+UX�h4ԡ՝��~\9^Q�W�Us�+�k���71Y �J�]r�W����8�h�jd�3U|������KUr<'��h�4�0UY��
ho�]qo	��N��J�zE��F��yR���|�y68����H���t�*I��'PAGM@s=B,ר�g�nN�nD��ǡ���]L�*���Ǒ�ct��_�;�~�� p-\ hZ�ã_�#�C��.�ݶ�6��e�VQ� ���͂�1	M�۶r#z'���'�} �}�1T�#��YY�������� <���;`���_"�i௡�@f�dD����>��'f�qV��I���

�WfU5��ԍ<���I&}]��8�~����$BPV9�t��p_%S|}�v���tR��v�s<Y%�������;��2�+��@i�7
�5�?���f���O�#�5��Xn?ȍc�Rn/�l�}�>W�<�.�"�U�c��}`��۲s�ߊҚ�4n<꾟yq������q�����?%"�<|'4ZVc/"�9����B�4�S��͉�]�c�ͨg�?z����H�Y���\�A�:ҳ.4�>��_��Zi�6��Z<������8[�N���N䇱��Q�)��I|���Q�7���F%ܨ������[�L�Z(��~�����`�@3pY��" �R["?Y�i^��"��]��s���y���tϦ�r�}�v{]6����jֳ��]�m����Qlw�?���]p���۳̫�KL:�g���v�	���+2�~c���T�R��h�PK   �rZ$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   �}rZ��@�/  �/  /   images/c6f01788-a49f-442a-a7cf-1585482f8cc6.png�/pЉPNG

   IHDR   d   p   ���   	pHYs  ~  ~����   tEXtSoftware www.inkscape.org��<  /IDATx��}��u��a����� �A0�)F1HbI�H3I%��-�N%��\W���]u���I.�w�h�mӒHST��� ��`s���g���3�3�0R|�C-f���_�����=_{��%�h@�%���A.2�D��.�"�K���A.2�D��.�"�A,r�-��@U>�h�~��(P�j��B�r�%�|`�C�u��:4�h6kN�B�lv�2�I��l�XC�(����3E�9�A����,����� E��k�=����|�T9�҈��8Tܰ�:f�Hgf2B$&�ۡ������O��T��^�c{W�NL&�|6��2�� <�L^f��F��v��l��������9'�4�ᴉ�{�8E�*�amN?�)ڼҟETT���C� X��F�߉�i�x�W����bg���,��f���$���i�X��x<m�X36w����5����+�AX��Y��uȀh��.�𓇧E��H�L��[-x�`�'R8D��KƉ0՝��;H�l�@�!�rC���"��h{��s���&�5ku+�+�CX��L��B+�$�����kzUm9�FdQ_׮
����p˅A�CN��xt�Y?y�b��ʳ{8��S�z�L�맒�{p�^q"�>Ofߡv6�R�˅�� ���븅*A�(��BC�WDrҸ�9��d�~Qh�V6���q@JpQ�R5(E�YʃI*VQ�b�;��MS�8ЈXP��Psn�	�/�5�VO����ߩ]�j��o��e�ZGe�N���@p|/�_��Z(8������5t�>��S?����X�`��݁T��p���q�ߠɪ>���~����ij�>\�q�����O�mDh�m`ⵞ~���^�
4�9�6|��#?C��n:U�������w��u�7s����'E�Q��ӗ}���P
f]�qA	�����ȿB��Į�a�]�_�����[�~��p�g�Z���y0D�I4�
o���h�^9����7z��=��T:�����/�ĒB�|�Z0�n^+W�4Wp$�2R��'��#��cj�;>�LpU]�ra9�o~]�݉��%�7k�ɚ4���>��ZQs��u©k0IN��������ʂ���˥ˠ&S9��Ǟdᅢ�é��q�����Z�<o�B"G���^�0Y:c�$���/b$kU8�a�əB��C�ɳ0�>��A�a�ND�0M�w�.��	��TS�a��w޲�{���4�Y��DϺv�aŊF����K���m%9] �iۦl�҃ɩ�y�r[R�8}yj_�ӌ�_�T*�g�?�p�|I�1[�n|����/�z
�12{g��&�~�#��#���;���'l�X��Y7~��]A�85�W��j)���\���C�L�d�f�1�
`�df����4ͼ���ŏ-��PE�!���#�|,
w���X4'�$�T,�3��=�J#�������3G��1S�q�p�	b�� ��}�Fa�M��j�al����'��<�*w�dE�L�`p$$\���m ��,f�gRxkoJDV��_	��,3��I���?�<��LƒI�'+�c���}���ӄi�v;cW��􎜘�Y��%�Wy�.�R��̻e�����c�g+6�`�"X!r��OV�����e�+�&뉿ON�k�U��r�n蹸XZ�9~Q��A�V������@�Ri'���^� �ALQ��|Q�	��p�0R�Q����i��e�vN87AX4(��m�`d�.��XS��q�UU��R�d�ᾛ��yMC�e�W�%�b�vbӽ��~�467��d�6_F��h��8�̌�si'�dx�0��ay�����[���`|�}d���g���>Y�#�;��c����G�G��8Z�="�בv�m��K��S�j?��٘���!6��\�D�f2볯�AyGF�}����=�������!�|I�X�N��N�U��M�j�nZ#>D�m���q�L�Q�3|��sx篒U7R�nzZ�i\�?0��3dZ����������ƻ�>����-lߦ�i]��c��hM�JK���g�u�q�'��B����fNbl냄��ey�s��-���;���b�É��Y�h߂�RX�K�"��k���\̢-�s�Be��Vq�j�Xi/8�Q�):�h/�M}s�ь���4��SL$�}|� ��P�]b��M@�ll5�!�9���{*�͊o)N�����ng�,>q��KK,��.�E	t�f�%G�%S���C>A��s��Wl�!�3�$~�"����0�ü����hB��3:k�pfm ^,����&'�����TU��K��p��f�Z�(XRiq|*m�;p�&��d��T��S,�ҟֻS�`A�9�pi�/~�tc���qlFw����X��kV9����W�󹯂�T�Ԫ��|��u�l��6$��E9G�14��ɰ�J���>GY�}.V���"�l�T�G>����J��|�τ��L�#s�s���#ٺ3k?�恗k2�ܲ�pq�UL�eXb��}J��X�-����|�u�ZL2OC1@�V1�z��(4,��#� B���͢�8����Mɼ�{*L����I4*��HL��(��x`{�:T[��K8f�p�tX��G��c�
�F��>z'�,:p�l,�*��	��Ń�]>ɂ��s8�TR�ln���/�y�NJ4��#b���U%8>b���G��F�r�q���v8$5c�x��J��j�J\�y\�Q	f�t'v9��)����+�����vCq��gpv` ^���
mN�dt�lV862�������a�U;��穘���C�,�|�"J[7oƦ�6hV�
�s
^��6��4V��᪍k��1Ib��C1
����p�
�b[��h����k\���t�=�q��p�'���rH%3������ۜP�̉#�N������W�"��Qr�r����,%Ϙ�����#1��3å�L�,#�;g��J��¨��Y(w&Ռ��/W��r�i�=!"���7pF����B�����9~|/Bg]�IJzn5�8�`��`M;��L���p��j��c���A}�` [�Tm�¥���qt2�4'��~'R���A��k�}0;��L�%\1t�Q���fh@����H,^�^�'R�n��]_nG:�P8�`��d8_�=Ob!(�#�LW�Y��x{�p���ű|o��!����^��O���1�����܊є���"N��A>��]�D�x�~���-�e�UkH�{	8W;����w��������.��Y�K[~|<?YZ����ڊD��l�g�u2w��ֹ��?����B�&�⣠�ಮ.Wr�oV�)���u|lz&IlN򵨠*/t�H�^jϜ�(��wf��1V���AF �nϓ|._[]O˟|.�U�/�$�d���!�iJ[E$^@�h�j��K 9���USpf�N$T�C"�겹�*'kJ?�������k��3� b׮]8x� 6n�/��s�M7��������7߄��a�^�G�l�,ޓO>	]�q��w���C�����{�ASS#^|�%��n=z��������?��^ۍS�Nɵ��2Ye?�s����@���as���/��]�Tw�W���F���t:e�\.lذ?�я������̙�X�v-�{�y�����7|���
zzV�	���oࡇ�f2S��3g�!n��#8~�#K��79���k<���,���>'׮X�}d����8q�.4Hp1m��U�5�(�-U�$���)���D�;��.$�6��g$����<S�3��1��s
����������z+2_9>99���F�&!�֭[q��!8�����Crc��jii�}���p�<�\s�������!�\Pѥ|cbY���8�47�m�땳�)y��1&'�9���恗��H֭~O�Y��x�1LQ�%��=L�r�����i�G�ƦM�e��?�χ|?��32�l����d=�ײ��P�={��_Ǘ��%�\ً�۷�9�Z�
;v����>+�\(���c��@i���Mn):N������g �:�T���8�\�4��זyK;X���%�g8�Y�������"�q���K;+g��/��;�C�?��O������z$	���[�A���9x�N�>�x ]]]8y���eN�F#��j�ݻ����E��u�]x饗p!A_I��0F�ǳ�9ܹ�Y���_
��a�7�����x���YTmq%��*�7�Hz�KZZ[���g�c�=�5k�H)�����|T>y�Y�3����|�+H&S��yvk�*%n��Iᐁ�!��?."���_q��Q�dǺ�	���kYt��:������L��W���#ô��yl���� �qH�,�ߧРX"��R|g�`I�����e���cǎ�ċ&�422R������̄�{(�*Ue��ה�e>gjjJڸO����e�U�Z0�\b�+��S�h�ϡaK�O|�Hڄ�T���q�X�wWh"� H�Xs:d���x��YԹP��
��^��V�Rf�z1�!�+��LMm�O�1���$����%K�ԙp�"[��FR��r��$�%+�|G��
z+�%��:n����t����ӋgBoی��qq+ �+«o�b�z�s�zf�l%�:�E�}��>�ϐX2��*\�.]�����	��}k�y���ly*����˺a%����[���
�bt�9���ŋ�g�yY��̓��,��,���Lۡp{u�%~G`|?R�����VCYI��L��dGw�4�%���sq8G�1x��G�'N#�yF�ʗ�)t�6��˻c�n�dM544H��l/�����ߝc���p�������}�?��:���(�O�fUV�_2���C��8�Y�,?ĲE3sFٜ-Gs�;.��)%�;�9����r#e\��a�8V�?�R�^���ͭ�:5<{2L֖�_ �=�s㰬�;�h�ae���%a�Y��g�b�!�J�o�?0�3��D\�v{�q�F�'V*����p
g�m�f3b$0����~R�4�qd<�]�c"�`1��ܿ�B��c<�����tև>�,�l�$�	Xy�+V�]U�R����� ���oŉCPZ�k����N���ޝH�[�P���/|��M� ��>�7�Dxr
;��ħ�S�"*�I�ܷ��/�?~ݫ��+�}H�9*e<�O=�^��s���_�4���Y��xc�a<�'h��������C����9=2�o�ݷ�9�x�Gq�έ(���P�H��_��������я� bd���	�|��[��?� t������G�`�a���-z$c��3T�J[X�M�ch$�[��)8�V��Ki}Dqʼ��8��:p������cV#����t���[Y��<���S�f�?��w�eF����z="e@�,6b�C��y�������{�&-?��߉�߼O~���`BK�I���Q:�h�5h��-�{��i�@�Ӯ����y��<|5<��ਠ�-��d�	�O�|i�����9"p*4�W�C�o�a׹9\Dȅk�u�V�"���]�K�6���^_�/βwym`t�5�$V��5�.�|�y{���ܻ�,ӎ`��*�E�F(��,Fh�J�<�2�f��e#Psw���c���&o��vr��&��A���9�+�j����q4�ñC��@���UUx�X��bJ_��M������
	��,�b^����E>�U8j����9�KK����b��B�?W���>�:ʒ�J�r�����T��^�^��_�Z8g���ͱ���"��p\._�����w�"��9M���׫�vI����N���&��P�
��YT��@^8��W�޻F���(�^?g9A��-�bf�9�\Vߛǐ	���)�s�Q"ʢ����@KG0�Б�u�> ��5;��"�����r8�j遊C�<Y6��҃;w��d��l{x:�������̼��	���r�b��3L��V�@��$_:�H��A3�6A��xy�1\}����?j��
6߰�D��6t��8���V<2�����������(���/s�c�~HQ�m�7��$i�U���lV
<�k
��1�X�����YxS��
p���
��y���h��X� 64�#��ĒH'R�"��'7�O8u]��
d�eMŅ �FY,�u���͋�� e;z��''y�L�J�L"��P�x�'Nj8;x�'��爫I�s��0�^��3-g�,�-��z��`��\Edqe։B�FDy�G"NL�t��!�و���xah1?Z��θ;p��I��Ys�cd�x\괬Ҋ�M�6I�c8.�U'�a� ����r�jطo����s��Q\�266.�4^�;w^Q��ũ�~ٺC'���+�\2�P�C����`Ȩ���P�oC�K���v��~:^�PK]��iBs�#O�����c���x�뿋-��p���s�o��{ﭜ3A�g�?�uS7�G�з���o���+�9"ԟ��W��ǉL:�D6�G��j��7��Hq1�8v*�G��]�������	x��]с������7��)�X�d������]v#�Ȫ��s����a<⦂�F�R/��v���m�hkm���d���hBgg�~����N
��я�n?b���t>���6�Rct"7O7p��z���Ds���/jey�<��� R��?Ě���O�����;�H7��X�-d��1|��&���z��B)6uaE�>��C��b����؅��:;��	KI�ps�8b149���)�r&ڻ.�w�D"����)k�=�đAf��o���F(�>gV�B���$\D�'L�f�Q ��Ŝ�-��u�&p�=��[9�E�sf+���F��"N�!�{���J}˖-��/�N%��U���N~���ۢK8?W?����K�x�wwwϻ�C�y����q�����;?�ή������]!��Šb�2�JN�^���*{�&�)�dg#�	�r�B@�Y`)��2��Ca��8��,����5a5�B2?4����ŀ�\>���-�΄�eK+i�[�������$[*f/��ޝ_i<� ~:r��~����u�)&�5�S0zb����l���(�������ʲ�����z�Y++GF�_%�:�:]x����������>��S�XY�E@N�.�p����ys'[Q\;�,U]���u"�Ek��q���T��gɬ6;�E돋l{K�l2��Q��T����q��hJ��ld�%��_�,�X�N5�_^1+4���y�W <C�,H�_$��7F��Rxe��S-r�p�a|&��<uD��yӄ�8[�X;,��ՃV��e���oD���3E�%�dB*h4=>���)���@A���<b��=�G������_��>�������9d�MȌ^�'O��a�TH�©�Ӳ��9~�+�^1�����Ξ8lQz�&���/)�|qy\������PNG�rVf����BM�c.�s�{Up��;��UD��3�eo J����P�#�e�<"�±8:SCx�<v�\|3ߋ�bˬ��s.���������Y<4�v�zxv���
d���΍��x�r�e��P���2p��(��?A��Y�3���yø��銕���kde�2w�<n
����$��q=5�鸆�g��}q�R@zrY�wU�H�f���beI��]=��LbD���M%)��_{=�?x#���Ѹs�1O�2���u~c�!o@��G�ᣔ �?)m�(5�O��Y���3�w�jpUqv�4L���|O�0ݝ�Eܑ���ԯ��M*� �?8~5YN8��H{:pV[�p�M:*z��a�/o�"��qb:��쥋etU�+�A�J��55��ź��o��,$]��A��!{��¥z��[t�]�H��-mA2��.�]��\��j��!�~�y$rԦ���R0��F8�8�AևX�/�C!cB��D}[�2p2鮍�4;T!����RҺ\�+x'
^V���v�ݞ��7��la��H�^քM������Y�@8��u�͞F���s5�0d��r�h��:O���TJG��6�XL�%K���])�I�L�/8�V��?���o6.��ӵ�W<��ǒH�,�Z}ǲЖ1<�\=�@���"�[f��b�X�mk�82�~�o�ɗx�������8�^�{
[>~?����[�.۵�t�Zx#�����1���-�ۉ�D�E���<u~�֧�������x�,���9M*/K;�.�]x��J��5�X
Xw����_��Υ/����&��K!o�+ˣ�-đ$��VW�Bx3D~��+{N���B���TӹV�'p��UJ�Z8I�xѿ(Q��h/���+����w�%C�:���%�.wr��Q�=�z�~���\|�#��wR��ԖO��������EVͩL3������	 p:�l"��DX���f�>�
g�Rmˉ�ŀg"[W#�h� qc�rٜ�)��n�A磇dD��$��o�V�U�>�����5)ܽ��Jp�S��އ���mx>څ�^�(8�%9�^2˂��H|8�Ҏ��U�.�Y���p��~�B�>r�x	ݱP�;��O��-��'vv������o"'}�.Gu�I�49�.����w(S@�(�B��(l����5q�J����IF���ɱhp�&.�,q'�ޛ�r����1����7шhM^R^^��]nI���X���Wojö.?�t�Dƾ��я�W���o�������VЯ�l�'76�S�m7���OϤ��ި|_�(L�S�}���uuN��p*]�3��x�d���Z�BA���>/>����)�f�t������HfY�o����&��v$5�ʹd��kf���v"j)�������]M���u(���b�������7wY��8K����|u�ւ<����;��xp�K^�G����jf1������d�I���ʶ~
�49�_�m���7���օ8�u������׶��v"��"g�MoW�4`c��pqSusʒQK)/6ζCTU2�0w\�҃Mm.�S������t�~��||]�bOdA�x~�ǃ���������K�ќ7>�.����=�Yp0X��ʎ ����xʋ�\,;���q�z�a���x��][]xx{�\���/�n���]W�n_���#��f]�7|�v�b�7��q��Z� �k����r:�`����>��#�d6_Y����,o#���q�::�	2��z�ܰҋxΔ��fw����C�ua�t�V�1�ݶ�K�C�Ů2�o����h��Fn�����M�S%��m�FȲ���v���^�d@��8P���,oi^<Q�(�@]���<���]6;ۼ�������b���Ek�u����:h�����m�
�ktH_s��_9�\f� �Xk�u{4��~v�]��E�������r�"��ŧ�Kw������V����٘���-zd9�b�Xe`�G�:�Qֆ��2���<D����5�Y�sїaB_�3�AT�F��e�4S�N��^�V��˫ZC��5�#A�Ө,G�*�p�u�HE�ir�K�d�n���χF�J9gA)Y ��G����d�z���?���y���2��;Ϥ�,	�,^`Q����IZ;�46#�Ԟ��Z��&jy#K�!�ҁ���,=�}X
��ұ�-T.3��7؂L<b_ˡs�*��z�v&�J��������R3���p��jX6AX�^Ff�C;:��䚼����C�xm &��3�4�%�4PƇax�aM�b˚4��Im��t�C.5�
b���9x�l�����i@s16Q%�x,ʞ���%�xyޢ����I��Kb`/Ze���/�`O�Oα�&X*�:sy�,�01��چߺ�Ϝ�o���]�������� ��� ���(y���2(��xq�D`j��.�jw�y��8��dӉ���r9��yrx��8��G�]�َ�p�9<p���+$�$�@�,� cΎ%����i'N �
 �0�t+��Սl&��iO�8��&�����\ml�o[���T�8��a�o��� ��/(�x�_�K��wb|_>�����9���+�'�K��� ��֝A���I�x𑇼��'��Uc+J���$��!I�\�T��U└�b{�mN{�}yV���͑�f=��C^4�� ӹE�;��A��r�e�1�[8���@�����8�I$t��%�>=�]�#;E0� J]�Z]z�/_׃�=?�N�S�����N�����)����x����.�/��VLN:�M&�zB������h�9���gs����K�O�0,��so͔]
�������	�H��rq����?/�Zxq̮�a�ۙ�P��1+�^����	���a�&�=��<\XU���#�w���ډ�f�\��T~�4���������7X��F"�����W�B\�� ��パ�p�m�}����u��q�e���˪I�W�k`+/����|MsKn\� ��|�l8�Q&w���D�l|����A���6?�=-���ɭ����A	;�J�A�u9xJ���x�>�h���p��a�-��$�z�y���<!���_��K�0^�#%��޸���h<��g����{�§�hpsl�;�e�LQ�d�8�j��u0�B�>[�w�:*I�/���{��b9Սu���I4T��ZhrQ�U�'l�9-o�t���tI���Ry�OJMtQ]�\A�Ӊ��_��	I���u���2����5r���j������:������<�Ǘ�Xha��健k���-�E�..Ҭzu�@�07��K�4T��v;ۋ�K�݅Ҁ�
a���S#;Υ���T����\��o�$�i�c��R-���&�^4��|��
��3G�	y��ǥP����I���%&x����9���kw�Ɠ�C���cx�Ė�b�>oW����ˇ?{u�V�s�Q�����`{K�nEB�<��FCY'~4���CY{��9������7��o�pcwA2d�ђ"�-ɓ�φT|���T.��-V��PAp��ݒ�('�����&�����#E&풞ʠ�iǢ�p__�l�WMBc�&y��Iz��YO��םR�� L�'�_%���?����Iy%O���]���r����3�L��Uӧ�S�䠅&WmD����\�3M�f���Xa.F0��}��'���y�jP@�G��JX81�+�3}����4�|���������+�^��n��ADH�xy*��2��;?���'-��<n�.`g��v���P�x������z�n���|D;��O���gc0�[:}�(�!N��WF��g���H"���[��y[.<��w6a�B��Rf]������D��,�d��FrX1s	��`���ź�	"��S���)��������,U��G�����Y�/d��KJ��o�uų������@QBH�+��*Xv!�\��7�8��Uz�\�&H�(��}�A��>R����O�\Y�j-�r8�e>oO�;?9+��g5;�Ln��0�oտ��]��^��P[�H=���{�6z�>+�^�A�]UDt�*�8�/��W#)DW)�e�+]���%��
A�3��K)��.��Fo���Y��q	70��I�r>�����	��d������s�1�E����JDʚ_��2��ˎ'{�L�9�͡�~�YZ��"�߅��vH�x��5"�?��S��e�\cUʖ��)bnXU�.��`�R���չ����,r��;�|���%    IEND�B`�PK   r}rZ���O!	 � /   images/cbf232a7-7072-4b1f-a35a-352dd9a3bcf3.png�UW]M׵�-wHpw�E������� ��������B�,���ݿa�=ժڜ�h�}\�fE*�I� �#~��EJ���d���'m6b������/H���/陸_�||HDT<2�;2�T����.��N�Wq�B}� 7����ˈ������f�?)a����禥m�ᣥF�K��D^���I���T�K�k����?���n��ZZIpۇ���j��Z6�u�F9r��'A��G����2�3�Ƿ��f��e����R_�W����O�?��D��O�?��D�������)q�Ӆ���;�"lkMYOc�c�ThM�� �t}�@+�Z[�m��U����� ����X�e:/3��a�!)���Tf-D4�}�h#7NJ�V��M�����OBT)r#��6�jx�u�u����i��B������$�E��@���n�������	
����[��ClM�m���H�)Q�'�SԹ�&h�B�t�v<?'����ɷ�$�c"�Ƒ����t���Z�;�h�ز�s�jL<a5������)�=�{�����F1g����l�+�5Dg��=�o	�w�^.2�P����l��/���+�9왷6�rZ�Q�L�e����$G������p̄8�8ox�7h��#!�/���^��ek�8�>�i����/�`�h,?�ۃ=�O��>�p@�$���a�_}NJ���:�����]v�s`��ёY����E�����$��"�a�k#�o.N�0u�����vm�Ǩ(D�����@᪲�����=��P0�9z[��#����V"���t�X���+%�%�a
�u�2�I��P�ھhf�*+څ����2.Uz A��Z�������m�1�����4g;�F�H~��Ä��NVV66�߳��+~��?:����K�c� ��ND���>����_���y	�0W�����d R�X��H�ƿr����,�����|��hj���^������יHKK;Sk�L���~�!!$���N�;�0��^��\2q�Y�^y�+Gr��:�M嫕No�� �����^�,��&C*�R�8o�B�z%�F9L���@�8��,���q���|=M�R��ba��Q7� �91��o��+�䪎@>��R�e�R#u�pU�<u�l"�)�\����w��3W7���l����I;+�_�(��<o��pq<b��=|��ʭ1�f߅V���Z��Ϗ�M��G�p�d���d)�yתX�����B�������/��3O"��i�^��w?iJ��� ��
�z�-�^'�����b<��x\�.�x�7�D
	{�?�}�U��0��[:\NU���f���4����fi����*���1[��~?i��c�=�̔�bw��fCCQC��7e��o�0d��貨hh9O���:w��L����u����d��d(�tt�,P��KȻ���@ p��d�&��P��<6>.��~��E���s�f�ns�&P�Q����B�?��U~��+�A��+�}R��Y�� e^q9eW^_?o�R?l���n�̨=`kZ������!���,]Hq�ʬ2�M��ؿ[�6��F$N���PW�X#�h+�(��`���R�O�n�ܯ��WV,8m�b@�� ���sfʽV�^��,uU�7���)�HR�磰��t�_�Gӑ��Ҳ:ĥ�
�h���!r����&�w�8�e=��o�vm�[X:���s��MH�s�Z�o<��sL�?J�����Ň�hۀ�v��i�z0�t��AKΊ�I�e��M6O��^���/�$��	���4G����<��4�Ќ����'����inW[����,>���τI�"���,olhq�~���xk�&����h\��H�f|r���t��DM*����_)��U�-dK��J�d.MB�T��W7p��dae�9�2s���KmZkZb���BCCA������UX��������.���h�����uA�>�r5�F[�Z��r��դ��Fv��/L��
IW��t�2l�:��Qb��.�6H�.{��3�Q�ވ���k�p�$���/�D.E�O|N��L<�©���l���!)^Z|���Hē2wu2r,.�ݘ�P��<�h�N�z����Mf�/\Gy��Լ��%y���6�h$W�K��Xm�E��>S�6�� at�W�@��oӎ���O�g{C�<\�MeY�o��x�l[�����
�zi)׹���)�K�D��ӡʌ�a#*.��T���/���
���a �ro�����C`|x��5^���� ���x����:!�j�֛��E .a�gA�0{�#Rs<$��*-��RvV6)��!&�-E���N�� 5�)�S�'��q��Ȓ
D`�g���Pb�A�[�As�h ��:w�:��~��9�������/��_��cO��e�]�r�Vr9��f����]���ᙼy�Cpƭ'q;�X�X��7�.�X���L�>��,����)^P;���ۆy��N8���	zw��f׏qSϭ��c��VH���!�"�i�%�#2��ri6kk�F�M�/f���5Mn�>��ب�b�О+�Y�	"CDF�>�n��p+��t*�"��Dx�ß�#Adk��W]0W���A�W^���u�䴜_�+"�Z���82ըZ؄E�z�n�C�۫��<�W�)�ni�]��O��~EH}��@X �����G�}��@��B��{�n����w"y U��-�پ��#+��!����W�x�2f\Gu|՞h��iמ���������}��˝����gWP;g����{r�٤(|�.[f�Ƿ�
ڲ�\E�ӓ�����uƈ�߮����>x���Tn��Y�&�Ѷ�-Fu�Z��	�U$ג�ݍ��Y�N2�/��n]��gW;��	ƥ�J��`%�5!�7]�W;��=#��.�M��
���7Q�v=��&�Z��0h�\b͕�\)��|<���)a(�����6v�K�'����so!�4�	���bŜ6����}_�V�g��9�d��ڗ�B~�_�i; �߳?ۗD���q�#�,TX��q�ō������665t���z�Е�Wwom�瓼X���/�/�WQWKk ���&�E��=<�IONOg�"'�+6,,��F#�����g5�d����;�s�e��Q�XN�6�W|�$�ڏ��_ǃS�#	x؎�9ӗ�zX3����b���}�"
ߓ
��>��u����h�y�#�ӎ�}�7���5ɚ2�jz%��g_��'7?\�����pf��t����2Ꮷ��格�Ev��&��1U�˚��i����U�
��}�:�T�����b �ς$ZX�'��?��U#ŗ�t�U۱㨎&0z*��9�g����E
±~���ZƇt�^Y���Xo����v1��!�DKMOQ����n	������8���ǙSu0�fbd�#�l�z�8�%��q|��^1�J E�p�f�D�n����mc����M*ˬ�B�W�ӎ����v3��d�ƥQ����{�i�����^#�We�;�
��>[;�<S�G��KG��)i8�D�u<<�K��w�=�����P���J�f�ǥf;=��?�&�M�D�Άd�lIďE߱sw~�����@F̘�"��i�,˫Uj���rm�(��'���T��QP�p(��m4�;�777���O�gl��S��x-Q�j�-!0�;B��V^��`B��eYMi��G��R-�oz��l&��]��t{\���OL��}��ou�:��L=Flތ�`2d���H�t�p�A�L�k��-Ϳw�����^nz3��:�g�>N�u�zc�7/�c�KNa�%�j�׶P��I�A�@rCNb,������X�-����1�_�Wx�6��=�����f�؈��\R�00Y��ۮ֝>��_�4��F�pe���^�0h?�>!/�=��R�7�wNQ���X0��R�ZQ�Em�"���E�܈�i���'�aCyƷds}�p����ߺ]7��'��K3�x]c�2������%z:�jk@Uy@��H4GڈƯP[/ �g���0�_)q�"���|�J����ٯ�P�ԁ�׎��X��٭��7{D�/g�K:���u�$�R���R�)?5�F��o�>;��_=uG������rЗYݯ�L�oǂ��>7�G���MUP?��`�U��[��V���s�]�KJ��z�O��(9���(PEx��~�I,���H)���+�߁�/��p��D��B���,��W]/�����8]ס�L�9�v�͊Ϥ8]�%��B���8J <�t֠����KKn��2U�
�v7Kccc#��0���e �e�n�V��wL���ù��M��S���X1��@��VvnH҅�]���$O��h���rw���h��N��򄜙�e y�2�)�8wr��]�~�`������E󦂪����4w��� ]6��k�=�>=��t}�<�'�5�c�m��͕���\�_�����P�X�QDWZ{ݽ�q^G��n~7���hN��C�S�l(&�.�����W8j��客6%�'<�æ$L��!�r����ˠ)��<��d�I���E�Z���7�bj�K�i��dI��B)��ozv�R��[�͘<�<�9Ω>��褶&�S�H����~��ʪ���޵]Y?\m�O�l��əm0��:�|���"��5jނBK..O��>�ҘR(����6�1_v�H!Uû��z
"�Ng1���m����_�O����g�/6�P]ʅap�͏�2l��N�旖�r�v.7��/�@v9O9�z���qGSG~��
�!!��4��@]����$��KY����ɓ�zZ�Z�����6�86�mb�-�鹭�-��2�.��к��/%��(w���6��W�/9{��ZA%_�L�����
�t�����՗�F���9�M0�h�/�U��l@��6��!~%'8I��uBy���j�$�Q+7�'�w@7��u}�\8�̫"҇�8����D���ں��©����n}�\�N ���8�t�L�78��U/�Un&�PJ�N�]�>p!��A�T�@᳜�ު��p�2HsƋ�Se��r�wM�qC�c�r-s����s��,.%��g'<
�t�:�1��_ط*�
�t؏�*���#���~~!5Q����0��[x��"ZsL��.R�r�]?kN�~�H��F�4�w�GƛX��[L;p��y��MGW����l���U����(��)?4&�p��b� :2���[\<����d���]4)i���?�>�/�WK���\:ѣ��g�a�UyƊ�J_����J2M���~�ILFF�/����)J�9;G���p�fm�ufJ���H���d�tquO;�¾Gqɇ�����[}��\�c��Mj�g����e8i��۩��
��kLz���z����K��Mw��څ�툡euuv	�nm��4[uN�"���/-g�v���Cj���g�ͬ?��w��c���V�\��|1j����0����~�_��0�_��L�Ym��Nkx�{'T����K����U�Y)�p;ɕ�����s4�f�;��]z��g�yҠ�r�Ԃ��y�����1[֥�=��ؿ�����dsI>N$�0q@?��8̅?
�$C�(���p	��WFj�������s.��1W�bB���Ŝ�c�1��'8�S���]K#I|�)���3�a�TjԬ��n�4+��bB5W
�3 ţ�1���z��{<&z*m�ԁ #��0v4�$���g;��_{-���e�6]��M�o��۞e��~�$;
�������Д��-����zw�z��Un����~�6�L%����U5�v��\�}��-P���g�H�8"L�au��VE�XQ[ۚ����$Qw[?;W���͆��'�<F_�^y_�4�hv�}�bn�A©�F����Q&?��N���G(H�?_�
O']Kg��_n�PO��#����}T�|�&���waM6��-���⶘�iy�3��>����(�vP�ՅV���dGCoP�R}3�<�jI�g�0�!Xh��x}��Jt6���+Ë�O��0���w���uж;�y���W��ϼ��m\s|�ّ���R�����M�%���O�Ɣ�;��a�����R��c/Z�����,�0�qǱ�~���X^������q�C�ቶ{�CIy��16�Ha�>�X����v�KZ�o��ҽ����3�t|��7a?��z=G����_�G������2}��{�v�1GI��������eW��V�c�/�]�{7D�|Je �CK���?ڠ�.�o���:n˅^V�mtk����#�y��
%�8b�芘��|�1�GN�#���y�sEc3�*[�9LU�b�FY ���2����5�5E$3�m���=��p��=	i�Q��*++WQ���e�@H�����\?;;���G%x��z���U��k��jX%|M����+�1�A�i|�W�wC%��y�k����z��)-=�X��1�6LvN�1�R�oa?��9H^��w�G�/M�&5����=P�ɍi
��$;���;%��'v��Zf.��n���d�	k`M'!����$D�v���|	�lO����~����Q�&�S�4���gm �Oe�w�NC���4�.����R��v��Mv�t�{�Ⱦ��(���J�Y�L��&�҅؏0����WɄ5�u���'	R�R��-�٘�,�縥�����,744���b�H��g�/�z�peќlbH��`Mz(p6�l�����������]��_�H�/��{���p��U��X?6��q�v��S�5V�NfR�T6�w�3=�����4����F����{�ZZ���f'{;/�4��<m�x;_�Q!�WǦo�ͨ��A-�W
��c��_
%��2�S���Þ+��D�Pӕ3�M*�����u4�����D�|�Ŀ�y~�e��z�i�d!XS?(����$��%�g�C'�]n<oI{�����^|�
�j9q��H˭f�Ș9�߂�U��v�rjѡ&B;���x��@N�������b��������I�l��1��g�R�j��rF;���{$��T�5k�6��C��_�oW����$�����U$�"��������e� `�06�`o;� ���\H�{P�`8u:[������s���?��,������$�g�4��r9鳨3CR+��Tg	ƨ���[�\��B[8�x�B]$�E,SE��{��y�����M�ϓ�T��zV"�Շ��\3�tQ���x���3��?�	6+�!3��׋���Z���*ZH�#��������ၓ��{b��m��J��_Rt���S��֣�Xʨ��Jg W�Ml������v?�q��]5f��w�5���>jzG��L�YE�D�_W����G�0��҆���|N��Yyu�@�&D/;�J����f��k_�$�_��^��.8���M��]G�{��d��9�1�������u:xK��+�;0k,����Bxn�.���Wr,�+���	mVjv������O�H���4�7g��J*�gk�)e�Lߤ���>�I>��[>�_���/[� l�B��A�qH�>a�mj%��^E9��V�<���- q:oyAQ�����=�t��F)F~���-(���n��u�݇�V���v�ƽ�Z����$qjS��ҵz���n��a���Ӝ�M�9t��{hv�*�y����͐���d8؏a���c[�* �
�h7ٰL�Ty����|g�D�CZ�q�%����'�'�N|B�V�Pyt3L2��bo�_ �R��O��1ș��ub��� w����A�-j;�`4���@���S����X�g�d�NM^<����E+)sNNQ=��N�`"C(h������-�^?[�b���(�>�|�VmPd��gUIU���h��A܎P�O�S-��G����/*k:��a����s��/�nVs��r�1_%�CҲ��P4��ĥ�?�@�Lع�}ȥ����F�.w��cI�7�3�n��3 �S�>�o=�U��������狙�K��Y:��c�����������������CF���0s�>�,�#��A����e8bD�����d�Q(��7d?o�}oA��t��}[c��g����g��,҇��cO�8��^^�#�<緩Y�_���c/��vt���OG��7�~w�*�:������ﲮΩ�rqq�0��_^����)�8�����N��6��-�nO�F� 9���\E3��mQ5�}���
�,c](!~��cSYN��/���f!)���2��>��O@��|S�
y��^��Le�\?p�vl�����a�2mᖏ`_[	�_XPJ�::�+��ѷ���!%�X<zM=Ȉ�]�kVK�|�tcw��
�j�=���	�F�N<B|v�b�e�&�M�����lؤ??;K���9��g�`gv������؛�~q��4�����K�Z.O�T�v����@Nf~�o�s)]�����:�����V�h[���@8��f�OZDDY^:�40���8��A)lS�ݘ8��O�VF.�F��;P����hx|�����b��l�(I��IYn�(C0�H��$��5ꮏ|ǈ�ț8��.="��a�S�s�Z��sR�!�S��ʗ2��^����h��������]�0�����*���-4�~3���i�E�+������+���k�Y�(�#
£i5<խ3����q7O���t�n��{tj�	��#K\�	)�X�Җ��H9�8e����M��l�T��,YR��TX�$���VS�z�D�m�{}B��m��M�9B���-n�ْ4����� 8������IN��Y�eVB�G���k��y���JQ[�G|�|n�/�ܽ��ra6W@k{�[�]j�xjq5"�A+K9���6',�ܭ��w�,A�1x���R���?ꗵ&�a����B���\���եw{��=�zn.�8* ?!TZ�}S��~_�� ��La�4ܐp@�[m�L-���޹)��plqU��0a?��ʴ�!�<8���.�)&��pW\���4Re�?&}�Rȅ�_�\��$QPy^��7iYk��$�Az��v�q\ x�[�]2���ҍv�I�P��O�G�!�n�77��;�<��e=RLm���C&T�W:�&·'�=�A`�[L��A��%P?z^Rͥ�q�,�Zxzy�Zk"c|��9���;�JK3�=�N����z���4�	�%��##�r[�q��n0�mv�3M$���u��vSc�UH��܅2�CZӑ��@�rr�T��ٱs��E2＾Z���$��yl<�>,X��"(0�)�;�s*tq��D�h��Q��i������s?
���A3J�1�ݩ�홢�l���ߝX�G�TB,�����g�WX�!;ϴ!H�s$Q�PF�f�Ec��G�B�Z%O���B�A.��pK�&�y{���j��>� �*>
�7��8��|�L����Ԗ��"�X˖��9'�8S����m��?�-_P��'S���D_�����Pĥ^�~W�������
�uXPV���F������X�J7E�'��R����y��r���n��9�q�U0�h_r�QqU�Ӂ����f��Ϋ@��'Nt���.��=�m��(�-�e1�0F6��PIS�s`��>��ʊ5K� �TE��4�}pa)����G�J��I�!���� ���d��&��0#uÛ�||�Y�%Mx�T�=���]��CJݧ`��r�h���p�A��x�4_���T�,t��1�Vy�(� {/�y��	,X�<9���4{���#cj��$t	��ڕ�_�bu���DX��ɣ��ץ�����4���m����8&�-��$�_EH��r���>^��X�����ɸ����h��$y����Gd�'iHx�[5}���L�0��Z�̷�{����L!6��f}��1���.3靌����N��Y�:��(z��Nb�X� �cO �_w�l����5�FD�yI����Y k����7�:�F;��x33�-v����b1���)20����3�q2#8�VG�1����_'М#���&��S&�I�5���~m�ێ������&k�G�T9ސ�B���e��8)Aß� ���H�'-0r��.�$oC�w����O��,��'��Bϳ�F_3�Ӧ}�t�Ȟ�iR*�P�
R0��x�q�q���1��y��o���^R#��=�M�`|k8��y��CRm)&Y��È��x� $"�0'
�?�9a�����N�c3K+��3�ӕ�/�>��6N U��JuYZ����}�<؋��c���ǩ�Lz���]���T{�'�Ұ��GO��&���-Ő=�f�h��-�~��}c�L*��64n���V8�H��Y�2����~I��DZj�%4v�M�:����L-��;�ED�7����B���D�@%n��Yu~I�;j� �8�戴^��H���]���͡�����䢜��q�/W��.��3+�'�U��z���I��ns�Td+�ڂ
>B8�T�SITT�q����'���{뉘�yO�95�Xs����$���Z�6�k�R䱝^8���K�n>F�I��L��wQx��ϲ�s�����q} ����B����x[��f�h��J��e@�N�ǵ�l���Sq�j[&!#9 ��|�����I�o�XY�@���I�#��v]fwr�ѫ�@�#�A�1b,rpp�>�b���1S<�)�?�w���	�x�Lds�3G0 �����{�,RqZ)�_~Ϫy��s:M04�H$a����ƥ���p1MQ���͓?�F�k�� G�f��#�P�Ǘd�bl�$[�:������M����#�h�x���X���V�����>�i*���(��� ]{��
��%�ma김ʡ���4���g����
����z�O)��1��w-H�_E��7�UBp;�GCz�w���N�L�0�5E��5�nA]D�X�ǽ���s;Q���>HB�Z���˯��H��$ik]�_�SZ��)h�I�;N�a�G����*f�w��M��IK.FoQBӚ�@��%�F1G�!:x:�Pz����⤻*ۍ��h���=��dCEE����}u�R3o|%0����5�{�'��u�E_VQ��2IH7��w��?�7G�������b�cY!�s;g���j4��}��6�Ŋ���#O�z��1�� 0��c�j�g4j�ש��zl�fc�Q˱�JC���F(�����V�{as榪�tͦ�m��-������!E�~rн����4)ɠk����9
=�/��U����^*���+�IZOC�,�[V�!�NID+)��cD��w5��4����%���&��$���lxk'K7��m\�{�qD����5T�%�9;(1���W��7�u�������Y�F��W13Tz/�B5kC��:���lꣻ�Se��й�x��5:���������##=bPGht�e�P�?"�]�ghhd�.:���%�&[����o�>�///��:*|���D�=����I����V��.��a���Y����۪i?]N63��e%�-����^"�U���eb_�?��I k�����@�@KCz�8A0�m�ܚ�տU4Ȓ��b6FqZܮm+�ҷ�8��z�7�wݤ�����p�� 9&|1�ߴ��8�����\�9�u6̀�v����z��?��6֙����>W㾮��}L�L�;J�ۛx#qoY�C������q|Z�>G�k �x0oP����\��?M����ISl\��/VORR,;��|�5�]��S�ω��K�5�ʠ�;
7J�)���kz���[�uY�>,���U�-�	�?4����`��z�\�����_�+��P��&�Z\4�dxEF���ń�`��z���/+)����Y���t�<;N��������e�BEϻ�~aɜ�OQT�,}UCWV�.�M_Jj�8AH�_y�o�,r+$C��9y$`@J���`��H>�*��ڻ��nV�*�*Vyۣ?��г�h���jUęK��}��E'�%fϏ�jc�rex?�J�/��=f�B�=:��q�&�#��E�I�F��fG�c�?��ή��"(�F:�ą��KJ�gdL����]]�ָmY��LZX��
����J����|S��Q[�r�����w+~�q�\�}ڈ��u��f;j�W������6-	���6�Yʯ�|�<l~1[�QO&s������n�t�mu2����ѥ��O���h�2��o�RD�);R��.��8�˖/!��f[��\ƙ�*SW.V��x�2�'�����-!w�ӁR#�9[ƾ}�����m�cED����#l|��'�'�&῾�"d\G�]lf��� 	�tj德����Ld���a�E��庢yWRa��٫��j��Z���T>��4��;2`�zn�N$ζ��C��P�xIfA&���0�H��m���*֒�uV�כ�DM�F����>͆��#KK�	t���8Dd&�qܠ;;�Y�^ M������8�W�1ݷI�azb���C�n�����J2Fa�l�s���Gg��:�t@U����w-�a�V@�q���=&�$esW��Ѐ))�kk�g걂#��s&T�il�y�H�ډ�T����!�/g��k�%C�!��hI�i�U��+~*|�������A�Ap*���X�^�+r��x��^ �)����!T++�{���2~���D��&����6�bC�n4��1ŚG__ێat���;X�_�:q�ry��*�߽q"��+�>c�7b�$wTJN�E0��2\@b��`;r`�'���4Z���i�tЇ�Ww�K��*Y�VXr����N$�j,A��7�d��G>�*RE��|{,���	4��?e+J��H�}ϳ����{�]W�f[J��E��U��q��Ӓ)�6���M�|��Y$C� &��S���;޺~��m�s�'��l"�b��[i�c�;��]։��HR���m��:B:l�;�`��%4��,��A��_��o�c~�Ѫ�ң�ŧz��G�޲.���kP;�^jbrk� -S :竮�C��#�☨�3�/`����Y�Y+�0%<F1m�,��h�pb�߈w�v�4���j�=����̌eH�HC���P��:� �α_�̢�W~C�����ٿ��T^/���Md�sp�^�� r#��5
�eq:y�R��kOj�3q՛Ms��%/�/���ө���\��"���s;(_�g�ڡ���]M���h������q����-���F���Qp��xp���YϚ9
A�)%���MČW7�<_�3ٚqzI}؊�z�8� (2����"�{��ńW��m���E�P�w��/5Q�����a����1D7�2mv��3���q��I�1c��Wl33sɒ���Y�tS
�j�[�<�2��W�!�͊�����Ơ 3j,'�I���m�7_Z��z�U�А�Dq7��TF��Ѣ[�����z3��kW~��X�&Sw��G@� �P�1.5^7�z�NSI��~�jlU��^C�TB�[r�$���K�����$�CN��ʸ��iaJ:cK��>�6�z�Ռ7��Sb������-�]H����$!�Yt晎m��v�q52�:��W+��T^��{F�u������>bw��:쭇�Gn�����6!蟕).ش��O��;?=�r��<E^k�j����2�|b���c��uO����4:V�1��kC���n��%4�2	����d/��a�7��a��ig��e;h�N}�!�O%7�o�#���;:��|�{�B�KC-]���iR\}�),�Զ���i��A8Wm�*�
���۸��)`�u���==�l X��fZG"lQ���f}D/�}��g���o#b�bF.3HJ�_|,,,���ЍX�ʶs���76�L3��/�O���j�n���c�db�		�@���"�l�0��In}ɽp�@r��Jƴ�����ʕa�SG�)�:��x� ,Z�ev ��q��LE�0r,&�g5��o��j�'�f��HH�K�{-ͻ��hY2�{޿?�i(�uu���I��Tx�q��1
9NG"d�c�O$D4ZЗ�^��co����������)ml���{xOk7#�@&C�P�}�$U2��%���eW���������n�k��<L���g[JU53 �������YJ�h�^P�ݤN�k���WsV�sެ��O�T�y�:u��S���=
��2�g�����F��mM%+��1�in�\ZQ���G=��ʕ��� V����U�6V���y8� u�>LQ0��!ZJ�3Wx��$DEJ���!�X;��p�#8.��bA1ct�~���z�O���������7����<�eA�N_c�l�r�w#���o;�t��ǵ�ϥ�H1����������/O�fᙓʬ��ErJ@%���ك���9ax�S��:���na��~�阷0bI<Rwq|(\��zU��8@O�Jb�+�Az���칻���khV-f�Dk����n���2�g�1��j��Tvm����y8���{�U-# �]���kC8qn(ÿՏ���OBu�h4m���mhr�-55�m̍�N92�0�Y���>�5�����j�\(C��ܜn��;�)�}㭈�op�e���~��&��&s;a�����ۢ��ltop.�%�R�يP���cƸ��ݯ��F�4j �I�U[Kk��F�U(n�R����c]T��V���_k8͑��T_cʑ���uVq?�{���+Z8Twܩ��"f�o}ꦄ�H��%����Q�Όn��M��n��,=�"�iE�6-�ZŅ�;�r���=Y��Ї57��ב��ZM8���34Ij�!���A:y`��vv��vh4,W�Һ9n��EI�B}��JRr'����bxyH@A���	�1��^U�mxV�g���D����̾��9�F�DF�y��2�M��\�߫�L?�}�'6�5��a\m�D�ϴ'�>�t���WN$�k���1�#]�A��CC�*�P��}�c��q�g^z���6ހ=5�F��sD8@?�6]��m�)���eV��bT�2`��.�b�yL�Q<C�@HH��C�
k�>�7~I���Ў��2����N�I���Y#�"�g�zY/U\�S8ʪ�\߬�LB��I:[s��}��4�-�����-GE���� �:��v��}�h��_~A�����(��P�=�.���A`\85�iި�����{���N�d�t�>I�>�\*�N�[T���m��,��(�4j���8��2V�z��#�����b��ڮ��>!�ԋT���Oˌ�"V!&8#+5ϭo��-�r�����VZZz������<+oW�Y�e�2�l*���8ǿ���<٘`AF�EKK�T������:�FA��W�P��s�.	����Z���8-�a��C��h�8� ��R84w�f���M?�^Y)��n�:���t�̣�y��©��Z[���ʎ�f��ݙԯ�0xDj����(-�	��
q{�;<6���{�&V7��6vB: ��~#��)R��S���PԨY��E�Fԯv�,��t�#�q��4r�tLr��#����1�z5�eFE<�}��
���H�G�C�Dw�Я�\�\�t%Ok������^~Z;�~-*��j����$/X���Lw�W���F�Z��������� ���6�g���B�	���$��?�@�d�����B���>��g5��Hw�h�p�]}�.�a��@�aēB2j%tg�/��r�� !�U�:_,o�b���$ǻ/���R�'�a>�t�xIvriq1W�(��8|�����ogi]������Fk�$��نà��x,�
��9�j"�N���E�j|u���:N�SeIUU�F���|���cu��Eg��	�s{x��h�a���+%"$<^j��S���9x4���x�D[(�F!Z�*<���X�4m�]����t��)���/_$~rX�My��N�o�8���i��]�<����^��z#'9GYQw��TD����j������Xr��&\㎸�TUU��WD�;Y��S�j��F�:���ʼO_Y�.'��J��O�Bu����[ ܜW��F�\@
�k��mǈ��\�S��	9����_���H�jQ�#$*��Lz=z��~GL��6����&�m�ݥKp������-$��]�-fW��s���_�8� =����uy�=c�hz9F�ϟ?V�=��e@��!����6��#����w�p�h3-��z�
e��a4�Xwʔ)���a[�+^'ЗW�vF�����N�B,��g����{Ău�2�^��C�"m���``�
^]_Vdᆨ�:�a崬�mI�������NtK(�u���Uq�L�ݑ����+:ރ�&n?St����-xa�S-9���a$c�q�I�Y�v�[Chvv0�=cW��]9!����F�_~��ܢϔ��2�d>��!ңzO����Ӱ&���C�I�q�;>�F3��|��fŊ��0m����g
F�pOww�U�̚�B�ݼbr�-[�M�7�v�nOo�7�����	�y� ��܏!ԩ�g./{�߈:v��O<�]��*�j�qڴi�����W^�3Q��NDNt����qL<5VGGg��7,hji�Z�K���6��'es۹瞻]�{dL�o��u���|�V�~,�i�Er��K���<�n�i_˚K.���^��=%�xxdT�k8���s;wO޵��]�v-�gK���k�<�.ǰ���N��C���)���F__�U_�#�y��)R����T'������ޞ����Ϭ�>}jG:��ڟ�c��>��ޝC�fJm�֑�I�L8 �M�t^ ���%�x �a�\�a<��>^o��Dc�Ѽ����tw�y���w�z��Zn�Ν��px�j�Je��qS�>��Y��&M�}��_�G�c^8�¡hNXR�OXU~��߫�p����3�4�Uz�D���&p�`4?��U���uש�*-/U�p��]�Ǎߤ�Rf����[n�X�'�xb>=�snA�j����[6�͛6k�^~��u�����3h�"VP�[�n=����]��Ӥq�6�?��A���;S���J.&�)�V�7e���j5������1ӦM�};V�q��X$=eT�;"�v?�3{����Sf��[V~�Y3���I�q+**�PK��^��p����F���-\d:�����1�@8>�a�-� �1��4�sf�sC,y�h�gUC�A���n0�4ۤ�nS������u��#����e������|}�e�T@O�3\K����с *��ΐ.,�j�v}u)H'���c����j�y�:��0\8TN�Sƍ΁z�E ��,:�����Jh�d��+�/uo����.�.v�EJ�y���.&�rg�^L��� t�`��!���U�5�7uӧ�O��^Vk-���F��kn���TO2�{����q����]hfϜ���poN�M�+
����I���5K�}��ѡǡ��r�)y\y��^�j�*S];U'c�~�Ѕ_=�FCc�����"�7���s}��q�H�g����a񅻔�Y���Z7�2QHZ}��a�^�p1h�B<84��R�P�q��[�ٿ���>r���Xtm_�PoiYܖ�yH6��~��뛚Z�M���s3X]5	a���{�[�(]�xɒ�����NXJ�,��?�z�����<��Ό��˽�2�.�а��+�$�,�rݴ���S��tP�.Qy��i��OJ;�����Ė��C�3��[����^-����w�Ɗ����LF�.ٺ�~�[����;]η���Bz�Y{hh(�aÆLOO������n)�=û�X��U�5���wɳjg[�[�M�����:�lٲ,��`H�%�UJ�i(x�A<�5�I������{��r�ҥ�R��;�֜!g4�x ?����m����V_��Ν;>����N��O������F$�|����/ڻw�E� /������w~X*�rnk�M����q�y��;�`ŀ���e��Y�j殌q],� �ɗ��e���'���J����6_��r���GT���U����ߙ�|�;&\}ꓟ2?��se�e�!��)�>�Yǂ�������~l5�A�9˾�⣡�\-���~���s��DCl�"TD������Bࢼ�'nߠ6Np?��«gUoinю�7�����@�:����>:hL���Pk\����7��H��K����|G���n$8&��q�����<��c�~�6]�sI����є9餓��{#",T�J�ń/\�`�Ԁ��v=�Lf<��S���t�x�u��̓�Ae-ⶤӐɍg'�>q}��u���D:WLz�Ld��p��k�f�Sw��B�m�T`ݴN�t\ ������X��#[�q�AWp���Xw��t/�����ZYݦh�	��WZ�
����
C�R��֯3����׼ƌfR���I�.�-�S#�����ɓ�3�m����g��0i�B��մ�y��dV�W���X4��\�r�C�vtt꾖,Ybn��V3o�|3(�Ǥ-�u
��=AG����(Σ����d���I[x߾�];�x>x.a^G�%�R9���b/�Ft���{��.�0|̞=�]+��L*E^zםw]��w_}@>[-?�!�l�U"D#���6:�p먮�B9���Q}��w������y���2֝r܋�=7g͚5��9�g���ҢǇNF,�ܽ��[o���k�}�C��5�@�R:j7�Y���D$���mLRU�堈���?���7&��O?ciC2شmGÛ7m�8���%��m\SX�1z��:Y%�yfcl�ʕ�\p��d2vƳ��#^xNֵ��YqF:zM{�c��.�	�rc�L��)y����?
)cS��(@���X�7n�~�����{/nx[���?>�`���9����N�sfԆB��h*�y�����;�UU]u�4��>��c�h�醏�����3{�;6j;�\����s���?^���v�4��np���C�ݷDdH��[�)�ދ��W�!�3�w�<��_�04����xEJ�9�.۝�Y����'?�I��-�N-/�\022z�@o�����w���37�4,�Q�(���3\.m��?���l�3�R.�[�__��Ư��W���¤em|,'L�������O�wU"�N���>v��~����,^\s�}��;����m��͹N�#��'��0y"�*jٔk���j���S��Os�6��u�U��ĉw��J���.$h�x�	s�)�萫�M��V�?��b�6�Q4�攥�h# ��X�N
���M�a��r�i�&3}�L�J�AE�UV:��p<خ��.��m�c����[������k�A��u��{�~����������^��]��"<7q����ҵ
Dx�(E6;�.k;���uq,�/ х�2��*D�:����'�H��Gؼ���t�:��L���&u��8�p�A>�FhA�����GMgw����}��i�jd�_�vS����΃���k�eZZ�LoO��3����8E]~ꩧ��/�T�����!n1,��}xug���u+E��D�c�C\Ӂ���d[�.%�	���N��r�e�u	���A�٤�^����<?[��\�l~m�5�[��q�ɨ��Fp���
3{�l$װ��_�f͚5���O�J:R�-Bت��)�h(*�b;��.:	����������ϟ5c�6�t����Vh�r;��ِ��/���~��m%����]~��o@D���=����vm/bN@:Ѓ��N:v}�yf߷(�,]�h���=�����}��n0V1���G<o�K��췿�ǚ>}�tB�X���C��Rƶ�)!9�y���Ү]<����f�N�N.>8�"�ہ��DC���Wnl��<���F�+��c�7o�_�x��e%��7��v��]�ޣ}����5{v��!:48d�s�<XOߴy�����o�{�[��������]5 T�<�?��a��k׮M�~�nihl�U&�l�r�C=�����w�lw&����-ǁ�VŪU��$��-"�*�P��f�[���S���Exݺ|��=��1Dù��e��혱~��O�8�R�nQbVeY���~��>i����o0�=*�� ��xMqw�>pagG�"�%��T�[6oi���;}ŕW�<00�,�eԃ ��{׮]	)���ۮ��Zw���T)���˿�7���C���������ׅKA>5n6���	�6���
��n�i�!�o�Z�T�:Q��tf:,G�#��גRimm�Y��ӕU�;��ݥ��}��O6��6�p���j ��1�m��5��о���������N�B�A�%�0�o���Z=�x�Ԭ]�V���y������F9T�eU C�b���g�q����h��I_��Ӈbb\a�aŊ��ѱ�C"du���F'	�}iQ��t��t�x�q|[����"|��[�B:)��i'�]V��eRֵ����Z6m]p��i�Y���ܑ���e�s"�y&
C�M��+<�M�Fkt�Q�O����GF���t�(��)5����:���Lʪ�tK��J��LʙO !+�Y���9�^��P��?��u����v�7���t{{��X�X��L�Zg�e�f,�L����4����c�`�6p�N�Q<�Rq���#,�<�t�[eEu��̛� ь�ߋBQ��ĩ7g�%F���3�C#�6&��~�z�ւ,X��wlר�	�z����&@�\ו���o�/��4h�X�����dQ�b1���pLh�D�,�Xv8�uB�pxF31�'&bLjfDQ4g(��b��HQ@�"��������{.~��w3�g����4��:~Tׯ�3_�|y�y��{���f�����2'�ǳ�<c�x�7�˿����k'�I��J�l6o�ƨ��X��g��?�=��O8�׿�����=�Z}/(<`������hپ}��t��j���T|^��ܼ���·����?�G��|�`t���y��ѱ��v��K_�ҿ�����};w,��I�[�۶ �-Ԇ=�����X�+"�=��S���_�q��V��3�++��Vo\<�?<|�ߴ���Z;��+��|��K��¼G=\kP N�+���Ɵ~�����co�w����k��F{��q�����[0�<�4~�$\�z5����}���k��X`�yu����'�����F;l�G%�÷���_?y��>������?�mv�S�Nt���W�_����y�w�?d�X���$�����o��������豣�e�-;���w��ݩ�N�..-2�1�g硏}�c�����C=��^�.�-�����»���W��ť�{-F���,N�?�"���;�7�m�u�B�N�M�g�Pi��]�Oy#��\�Q�����Tj.�H�����կ��y��>h����+v�\1gΜ��-<���H#����9u����� � k�v���>�/͇?�3;=M������������̿Gi�_����b�����X�w��M�Բ���+$��d�\�z�ϧ>�I�jE;}����y�b� �{��u�m��u?��7�w_~�đ�E�A*�� �C(w�*d��B�m��wM��
�zUSS��2���*<��8'y�b�R���ʜ$>&�{-�j����o}q�J��!|��ʒ9z��`��n�ͱJ��"`����@8 }$�4�)Q�o�h�%����P�������z�+��Ϸ���F0���	fdߓ0~��t�u�n�X`��B��k����/x�~�'�9�< ���c>;=#���-3oA'J`_���������w��>��ɼ�m{��&�I����{�����7L����b����_��" �ɠ������6K�s�M��KWͧ���T�A���f,X�PJ����$��G���:^��@a{�<AދZ��?�ն���Y�_�U�����6��ѿ6��ۿm>�ٿ O~^���%q��v�U�U�?��gM����`��p}��uec���b�k�n!��������ڹ���t�%����C�������ڹ}֜;{�\�{ `(f �}h���R$�/l"WS�S�P��
��Q�fa�����|��w���o�O�����v���v`_�¡!���tK���j[��Ǩ1T�E⾹r���SO=����c�3<��E���͖�կ~���`����s;���V�A���k@�ԧ>�ܵs��{�}�<�s�d�P�+'�=}�����}��]�v}{�޽��?��7�}���NL4W��-q�JI8�����\������/�������6R_���췾�����a��� ���/$>����?��?��������a�Ν;�}�ӟ�gT�����ʖ��/|�<�wj#��tٶ�ѱ�/~�U��T,p��<'h*�Ʋ���ʩtrY��I�g�s	g.
^ ,���aђp-�1�3C��l"�Cy�P��Q�ΐ��J}(�+�'ᵁ�c}��Er�%�������_�%&*�8m^j���E�T܍(	�{�vM�/x��E�y���!�1{�@����c���*Z����jk������I�&���o�Z�B�o(�0�,Ďs)�}'���u�5�Ǥ��+�xB��V�2�,�2��r�h o�4Cʳ��i���X��doؼ��� ���>LN� 5�����[�64Ւt��y�㫅��3 0���vS�Ke�`��U�%J����C�V(���<���¦�g�1'^{-Wx$Y��ļ��`����9}�,e �E��, pP���6���ٳ�t�g����2�N�_�kMې��ߚ�p�_Gu�s��{�D�@�E�X;����̪��>����79����7�b������)����?��ghG��E�H��EyD���~�nas9���%��`���&� |�U�J�=�� �z����S'y,�e �x���G������sO���b;]���:A �z�p��>}�o�;�y��>����B�c6��~<��������F^4��j������o|�}�++>A�1��[c��8����g��5w=J��)k�~f��~�g�j&=���Ϛ'�񤙝�5g��_|�%�����.�0�0�H����O������������+�����|�{�.$����jܡ�c��ѕ+W�?��'ãw�=��C����珛��s�.W���(���R��'0�w��~�|��/�_��_� ���/ Ø���p.�_)����z?�p�g>������{ނ��f���,�Zd��[� �En,�OC; "��sխ�ch.�L���b��(}'/<�b�8u�4*�z�����p v�M$�,��bLz�����y�z�'N|�j#���C��;w���2�	�Jԡh¸�F����jCcs�g��������q{n�_��k�0�������-J٭װ�e֐	��f:��$d�y\%?Jߕ���	���ʹ�p
H�`���zH78N�yM\� q���6�2��Jh���1�����t�?0��7|3X=Q�;�H��f.�{� ��n�:��8 �q}D
�Cm�N�[d��.��;����o��y�+_��+�"��w��W����k?��j���K�4���dDx���u�,a�o+^x.w��K��{�<x��S�����XfK�,�t�����sl�q|u����g�2�%`מ=,s���|F���v�����X�?EѠB������3�Sػg/=��F��@Xe�(� ��y�hd��G�����g�%�Jhii�iO�z�]G�
c�� ���O �k�����$��u���=���@��w�ޟj��u�N:�&�j�W��?f��ܹs�ݽ�������8��C7O�055K��ŋ�|������"?+�I3`p�Zj.�����������_��P a%@٠��%8�� ���7��Fh�����$Z�X���12&�SQ	�;y�yᅗh ��կ�煅J�}b{)O��8z�=�hX��ן$�p�a��u#)}l�|����/��5�����'>A`<R��.9�w�(��h�Ӊ�-��饋3���i��Ëq�wׁ] _��P-b��P��J���K)r!�5��$�ј��M;���&5���I�T�L8·�`@�螻�e����+�iqjɊ��Ë�zcT*�� W14z��1�eLq�]�jNڹ~eY�@�f�r��4�O�$�m�����$Lxq�"�  ����EEt�����"�}�MKek"�5��5M��w��6���x|���L�Jzݽ�ݎ��Ԥ�4�e��߁�I[hJi��\��A�^;{N�W����y~�~�Y��a^�6��v�;��F�?��z��+���N�2���	E:���������
����`�RFR�|dɅ�����II���Q]�����N1b�Np\�;�����g�v	��ߵk�����v�b���{��kn�������R�-<�H�l����0�`_h;N��n���A�̊��R'��p��; ģ+�l�Ռ�kkY �nܓd�˗/y�?�������}���=�{p�`��ˋ�Y���n��xo��ޭ�v�x�,��W^y���͂����C���0Ď�JO�{���- Bp����z�`���W]ZZ1��w�e!#��	`SB�!:Jϴ)�m��O�O|��(���� �GGǝ���K4fK�!D)ܯ}�k�����<���ͧ�e���wzX��%+�v��ɟx��7�i��a�qx���1A���Th^��������Q��G>�s��Z�Qn
�����7���>(;��.oX�3�8&��P�
�x�e��~�b�-��lP�]�#����8.�eR/r�뉇0�g�V�m �oTܴ\��`Z��[�x�9r�Q��腲׃��Hy�{�o���G���*A��̔��s�O�G�!ah�"��n�%�\B1x�����ΟvV��e(I��9� >0gEݠ�pP��X������oS����3?��N��������3��s��k!��*�8��)����y��oa�N���w�ӗU���,t�-;oQ�$�W��5*,L��1QP�c_6Xq�RPV}H��T�c��7��>��A@V�1���
h���-�?�,r�S&L"Z�H$1�^Bo.���᳁y*�s�������r#@K[[��������v���+/�j����͕�W3�"�NPQ%-���s@S�7�.�;�<hN�c�{��7��?g�sX<�������N�I]
2�<��(�W�B0JG�AbҚ�K�^.�����F���������`����b�>nm/�8�.\���՚Y�_0ϝ�>�����vތ��A�x�a����i��1���]��"��a�&��ˈ@��ؤB�FK�9���E��{��r�t٨�Z��6�k�/��H9��J;�̿��23=��G�ѧ�35�/�$�-��ݶ �-����݅��.��]4�_�~�5�X
��Nc�J�*��<)�Vl��<"k#��b�;]x(�G �3Ky����I�;�l����E�tba�`���#���0�L��F�Z���1g�ޙ��X�������l
��IV����5#��g�#��%����[�EN+ Bh�C��IXҧ�16m�57�4���!� `R�X}/�-���"Ii�_:NY�VK~GB6q�gB�Ѭ~Wy������G��^t��=��s�X@������{-X<>���P���o��y����$t��xM���6��ҥ��햄�q�W�\�b77�}&g/ѹ�8����8 ��'zC����奈�� �#?K*�B�
D�$s	@t 7O�xʓ��]�|1=f% ����YL���e���?�7�j����q����s�b���.-Ų�޺�dV($�\�P���,�����%��|S���a��}�s|��p����7^�F~�NQ-YX^2{v�!H,/�D���<���OX������/����^��Պ�妪)��F��t�B#p M�g������k]n�ґP��)�}��g��g�t$���H���t�["2� �������x��]s:ߐ��#�=�;�m�>�*~�o�U��t��=�o��x"�ؠw�~0�
���'x�U3��e�ӟ��?y�#�xtvfv �s)����߶ �-܊����1׏?���y�[ �0�U����	`�KP`�&f���.�ˆFꀗ
��K}xx�ࡂ�w�����gU�`_�Db#6/�J�{13��)�be�I�2���BP86�#�(�^���XJ4��� ]�N�/dX�P)�����b�`$Ո�� ��b�HV>8�m��04�8��a��)
x�,��=K\N�w5ш^"$Z�p>ME�.������66>F���!u��>@� �Ÿ��Y�Y��&q�<��滯|O<���+-x8d\���e>�WX0S/� �!QY��<�B�&�c�<�lQ��؊��b��>AD�N
Ev��O�!�Fi0���I9��[��'}Fֹ��=�^���E�˿�T��ʀ���3=V�c�U����!݌2��Ix����c���ax���!/F�t�9��#���~�@���oG�*y�CG3��>�
���x��k��k+%s����ٳg�T>K�j/��p�J@�>�S\O?��x�;j�6��,�h��u�.�I�0�)�����l�p��v@>��ʲ�H�TI?D��S���5i�O U4ȼ��3�&�Ixh�e�Lr^���9WZ���b|��&@9Βɻ]�N�Fx���^f��Z-^�� ^����<�_|͎��[Ϯ'�![�U�ߓ�	���Fn��?����7����#�^��[@��/m��Z_��,��.]���:u�7,(� _<!+��Ef1E�'bN�2f��8�S�[���3#̕Bu|)���g�CC(ni�鲂-�u<�����?p�`��k��7<L�����Z�	��������<	�3$٠�x^�֮�Ð�3ҏ\	P�
�8��G
)��} ߳���K���{�1�aO�,��aD�?=�ʹ�-Fj֤��2p�+<� �0����w�|ZZ��}�M2@��K�?�b�}��8j�3�CI0�!y��>x��[�e<9����gժ�MB�Xe�積��O�Gг`n��ҫ�p�}�&������ �Y㙕E��-Z�� Eb �:�����jrp+ h8�e�J`�EQ
)�k%!�P9�a��Gx�T���jo��<���Z������v'����$�f��zR�pm��Ŵ)�m��ĦǕD+�}թ��%y`G���eDS|n0B;������tC^}l�WX�r�n�#�]��JxA���u�#G��b$TM�|	�#$/�Ɇ�6K5׳��$ɑ:V8�(�D��*����T�P���������r��`�FU`�l=�oH�F����{ *���Q3��Hy�}�s0�r&�X3��q���*C�Y�h�R��T/^&W�k��5��2궯=&�N�=Yw* ��/|�������?���;�u�m�ۿm�[��0)%;�n�=����xp�����	s͂I��+�n7-P
kf�s�q�wx"�U��`fz���\yS���ӑ��F��0�QL�/Uw�#_mZ U�ɪxJ�0��5�}����]4$��T"<;��jR %sl����W���%�+�������B璋L,�?̰v�B�5�ۦg�h�z�T�A���0��_��� ]Ԫ5��߱�	*@`a�uɢ����;�P�* -fiX�-Г�B�j��;Ɔ��+ٮ�V�\�f&����<��o��~� �7�|��{�f�1���������r��j_��|cqZ�C�q��P�g=���@���]��v�������<1w*�(�t��. ��!�zMx��f�	o�n���^����,����S��0li	���k��X8Ѕ��Өl��������R*��sɁ����?8������K�����u�L��LSo-��uz��b<9��3�s����ת,�W��խ�7s=��!��{V����zΫ9P���f�d�R���pjC������r�Ŧ	X����y�ǗDa��:�
����7 ���[����O^-L�����)2f�8��?K��u#x�2�Ac���F�bm@���$J��#_���m�� ��H�a>�E]=�^�@<�G�>j��?������,�L�#҂u�p�|l�rc&E�~8z�Z�2 q���ȳ\����{ߎ}����q2�6��lF�')�S�M(VQ�#������(m�9"���\�����Wn�v��t���'��N�KiF�Y�y��z�q���1��97q�Z 
���'��$ֻ�5΂UW��;ne4D��C)��(�{�L �:����KW������������dvv:�M���y�ݾm�ނM����gw�ۂ��а�Q�M���������3��x:����{Ԣ
*ݢ<��}u@O���i�|��Z�:� � 5I�[V��8]�'R��v=�<ʉ���~��=)"��UML�6�X�U_ ��Iɨ�/*F�/�:��<7��,؆���5�zo����4�'M�������!�!�A�D$� {����&-�����˂"
jn� �r��uȄ8U�@�X	�����'��f��H\{�yx��A�YmIA�@U2�O�y��[jJ�����1ϲ�$|J�f����xpK�'7�^��τ���@2g��D$�T�L�φ^v�-�|zd��<kٱSDI
���|��+�<	vA{R��,&�A?ۋS�b|��JҘF>��0�v4�l�y��(L�m4hK�0��w��zp��x�$��Eހ�w�u`�c����)z0���T�8���W��8yFҴ@s�����zQ-B�sSF���u� ��s�WM���-��5��̿��:E��tn�ZJ���ք<��
_^�h���:�=�ꌀ݀No�xΚ��UI�9�~G,w����+W�k{�>>595�DH8�-Ht[���{�5���Պb1�)�%.�ϝ;�߮��zP5�K��M����&P�J �!=$)�w�Ŭ夐Q�z����!0���QT�Bfn`d����4_5!鍬d���,;���MD[���ȫ!{��jj�`HƗ!tj�F&	+y�����"��z���0��z���=��~�#�g��_�p!gR�s+(�AO�5�\-� ��eH�xh��-�E�72;�������Qq0�f6	?����������S���%��
�Z�����D���E�`���ؠ�XܜNj��_���� bޔb�!�1�Y�>Fq?��x��<g��(����Ɓ����3��+ٻ���s�%��J ��|�J^�iO5|��Rw}L�@y3�j�e�q�rml����_�ʧY���3;М!��#M	nA�R��ӓR��~g��_y�%��NW�5�K$�7I��{!T�����h&Z�,� �nǌ����+BCc!D�>
�a�pM
l�%�&�n�4!�uI�YĦ�;ɶ6������
��hR�^�i��>��Ŵ���D�4�Lij�P��R�Z
m`so. -5���s-�X��K��1{�	�!��믿���^�[���AXM��l�ۻm��[���ֲ��++��?~���f�BDq�d`�4 ^��{1�4��
��јL�|�ܑ�:+�V�����Rr.��J�:��D���,�s�t��6�0���"��E�8o�ϸ��N���J�!�2�8~ʢ� ����q����U� )�
��1�^^���x���l��i�I�",
�%B�:�3��H3�r�2=hni9z�>�B�m�'X� R�� Jǈw,U�yA�]@B�T(0�I�'</۷O�qգ�����&/m��Ԟ��Ao�z9�������7v��~��lr��R�o��0 ��b�bXSp��:��+MCq�b�9ߔJ��Av�e�g3��3�'/ί�6�8��kT�P��F�w>)>�! �2Y��4���͘��C����W�j^;�?�b?�)��٬�ݠ5p�'�.w���k�Q�@xf㘔<_J��q�g�T��<)*T#�Uc h�徨J��G$�}��c�����X��J��-6�~?�	x� �8~�"�I��NF}Ძ&����=S/%�*�L�(�B�*�Y�N����PS����<�_<�ӏ��zc�;�zo�uwo��:ޞ3���k����� �П%'5�J"@�����n72c�U��b��x!9L�+�
� }E&��&��6}L>�$K6 �!I]�HV���-?������+�J�4xe�����9#z���
J��V1<��0e��T�Ъ��B� �a�(�"�/�7���4���h�.G�Y2.�4�~�S�N���e(�z��A������"f��Y������762NO�/�/�C�k�nJ�l߾���]�>B�j#��f���Z���YV�C(�ew[�1J�M��9�� @��Нn�S����Q7�G��Պ�A\ނ|D!�qC_"j��1�RД���(�yԼ/�"Skƻ]�/^Y(t`ަk=��1+���R�R���_�",ь�M��eP_��f�ւ`}p�|�M�kt:�^/+�e<$�Vh��#�j�j��؅&W|/�2���>�-��A�cρXn������c��o~��m�=G�*����V��Z�N?�u�}Vk��G�1w�u���SO>M�oآ��wpSۨ�r�C�\<�N{��o�:��k/j����U��C�l�Us`IpW�HI)R��0� �t���d��u �Jy^z��|	PkmvI�.�V�/��O���bbl��H�[����Dn��*�_�f|�l|G4�c-t�&|y��q�%�G� � J��*�xrMS~�S�Al���g�-��^z�Е���n��=��Λ�s����ཅ<*�Vwrnn�C ~ _Z�\W��b��F�/�?x��n'L�'�4VԪT0S\$c��p�\����4�)+�/j�s�s�9Qi1b�Հ�WBdKN*��=&8�j&�3�).�xbhYh9�C���H�c�!s�aT�`���W����[8�\���]�M�)�
ͦ���ga���w̸������2�@l��5{��1�s��J �+xc��h���ǹ𹸤2��bR�A��')ñ�&�d�Ɋ	eetb��j�
Oa��M�J�ܯd�-}�xґ+j�[T1�8﵂u��MJ ��I�\ҕ<%�Byd1S�. A+s�7�W
^1���Ɏmԗ4��oz�r�T1䞅�}�R%n~���6A�7�6y��8���uC�p�\�� BCR�*�ȈƷ�� s���b2�+��+h���\ d1�9�*��K�滯�bN�:ev��i:�v���H6Ҡ/A�&I��p(�u���{jӒ�9��0R췖Ne�e���~>�yh ��`Ӧ�^<�p|�����w9������u�-�d��8�z�Ai��_�J%M��������s�*��%7��U'
���~���z�7w����Cwy���m������>7����#���(���XC�綟����$�������1�&�߅��2D���^FC��Q�S��Ja��4�)J��Y��Zp����.X'��;�Qq1)�fy�@>�g���rh��:aw_-��	m
�e��������[�h��%j��f�%��Xc�V�Ux��E��Wh־�$B�Z+8W0��V��W�뗓���zK7S:��:=]M�Ӆ��$��.�ߘ���⌦�ϙ��J9 v�ȁ�Qʋ��z�����Kz��Қ}zs�5��o imö	`�P�mr���W7�h��y�� �i���%�wî�H�	
RwYa����,6H�h�+O>�O�?��ˍI�P; ��!�M=|��f�췾�-������4H�����b�C�[ ��x��P�e��W z��
D�ɦZ��
�FW���� ̊o��E�����Z��h�|���Q��wk���X��K��	�
=�By�r���O|4�/�9*�J���4�]r���&!�Gu{M��,-.e��K�ة�1DI�9�˗_~��>����8}��o�[�m�[�)��Ϳp��אַ���	�n�	mѭU��_qU���fa��F]"C�lG]lS.` ""����^�/��ӌ校@-b����[��^\�	��X�Usz���/�C�NgU_A�o��i�ɔ�qQ���$	���5�u	 J@���d.��LnN-A<�~F��DT�B�}G�B��uy�U�`�w���,�S���"&4��S=����"EP�P�4�7	�ϛH&�(YMU;��ܩz�)_o�ë��Ip�X���9�E��E4*z{A
�R�$� �..6(N��֬�Kŧboc�o!���[,����OֿJ���e���^���a4�5�Y�{����yS{!�XK�P�@d ���Aov>��چ�?p�uS]����$�b��x-ziT�k�+^o���-S~p>�w�(��k��y>!G�v�����
��w(7hb�z*�[��^�۫�t#J���z�~���u�9 �<TQ�̶���*�_�ח\	nL+���V;�w��w� �0�$;�����H���˫�,7�9&t��
~gE9�_6�Eo�&�7pGD�B�l\���þ7�}����j�u���PK�r���urii�]ZL��ՠȀ��e�-!Gx`Q��4S���ٝ/C�Q�$����M3^f*v�ﲞ�x ��E7��Aۑ��e�R����ݔJ=�'�)�+Eή�Ŝ�:&�����H=�xb?�dTn�X`E�>Q�����u����ȅ�K�Q�g�9���_�Wl n}�eiu�Frll����Q���\(J$��9q%��āMpM�PD�ڐ�G�oVM��XTR�����Œ"����:gΜ<c�W�:iA�r&�F�eN�%?��;l�gN7��P��ԏk�X*,����h(�t�(�䅨����{�S�W
�ę^2U��/�۽���bU?{/���Q���L���  ��q���Bѻ��rv!u�J�ٿ;���,(J`�yJ�� �v�C�Y(_�B�q<0�#W(CB�2��;�g�T6%�J*8�rjg�s*�5y/n&���yͅM�&\B���׾�B��GU�G�Nƪ9�=��ɊBM��E�Nnn������G�{fS���w
 n>�q���{����Q�����Ȉ�sǎ��у��<�a��.}�4�j��U��9�%�:��b8�":H�^N�q�Q�����%c(��=&����ζb~�����n��I�5Z.JrU��:?�����l��.1ޅt�R7#��0�v�)?a�'F'�<l1w��xȰA�Q;?�P�B�=l��k6�m33����i391mמyjBs<aO|/�t�����ٺBGL%�����Q�/�Z����u��cwh�c�3|��x�ڵ�����vcΡ�ΧT�4���^�("<�nCR[ZZ�۞�����n���xo��S���+��!Q�$@�E(��UJ�ӌ�[�d��l�,�ѡ�݂���Lxp���~6/{���˾N\�;�L&���_�VR�
�����v�rۨ�W�EϨ&|d^�RhQB�iC�/o��U�j����JH��@�)a��=��Y��gzr�t�������k�
v�@(�/�o*�u��u�?�(��/xzr=K8E�Hɜ�G6�f�JP��(�d�p��1�n^�0}�ϕC�H�5���]�����Q��{��:o���M�3 �T�䥚��(�2"�s�[P�PH>�&�r�:�A�j�+�"07�x������=ٜEYāIGAž�0��v�vї��t:��f��N��G�>w���UpAIY���{���Dv��Y���3~�]����x��<��򀭏�@4r4���̰����d���%G1�$��Q�����z.�j�L��W1y�צs���7O�|ƥT�pj#��hZI_�8�g��}���?�fD;X���7Z�A��\Cq��P��3��׷����|ZhH"fI~�h��F]��H^��Eؠ�6��4*�sQ�җ�B��M�x��ܓ�t�]q!��˿��C�}�l�ۺm�[���m���������LRk��3E�2�&%�S���q�5D:GB�����x���Z=�Gd��˸WOl�;&�k���4Z3N��J�k��W��j�"@�[�v��N�}8��W�qu�k�~��T�_1���{�-����!�[�5ʪF:�'��5�]�r@ 9��L�5�MH�l�(� E�t7��`�n.Z��fM��P��f�4��\k��=�¢=W�ш��<����e���qN#ɤ�Jں��(ݓ�J�F��)�Zձ;6��>�vvSY������-����.���:I�񳍠o7�@��=�ݾQ]g\�Dq|��C�c6�<�߇k�=�h�{P�d!x���`j�RȌ�t��+[?�W�sY �������A�!�f2I��D�U8� ���%z������)�O,���M ���~��[��si@5��J=ΈJa����F���?��Re�5�t���רpL�u���<o뵌���w�YS��*4uWfX7���]�*�0���E���r�#��x �Kt2e�9<����m��.�~���~�ҝS����_��G���M����>[�o[��m����6�n��Kms�e�
}���s4������e�Me�8p��B���Ё�A^��: �5��KY�X|�b�Ut���B�O�����2�Ϣr����7{@�^��r�Z��"MA5��.�_�	(ȫ�Ui��\���F$�8�%p�N��K�HaI?�'ޅ�WL%[��FU�F��L��B�Nn"�4Y��YE2�)�6:�ysu|��L�s��<�(ƀ�EQ�!�4���fI{<��yu?_,�:�D���+��V�n(<� �	}��!\Ͱ/�e$e��r~�W��|v�NWHE<]�v�r���T���(��W����@(���pE�M�w�~�R��Q�tί���������&�1��ތҐ�:��);�v�7�&Ѣ�2�-F��O��-{^�ZH��)<������"W6<��mJV�����H+���{743�?z�:��� ~~#ٹaM�_��Fl���z���%�#_~�6%��b͢����j�sR7|S�6��r�Q5��7K��������d7G�ɓ�bS�L�[��!vJ1
�_{����Vk��f�ݶm�ނ���գ�ϟDlu���Ԍ��6��QCnX�-����hi��iiڑZ�a���$9�#�S���8դ��-v�.�:t@E@X2tA�Pga")-�#���j�JΧq�.1f�u���H��B��6/��^1F�4�k�e��rg�X����(̐���<ѫ�`�>���0Ι=u7�5֟�̀G���Z�t^ߍY�J���ȸ� ׬jZ-�F�,���}�̄�����kxYSѨ��r��/�(��3PbXCo( �^�,l�iyV#��`�\��"��"PD��hqe���P`��xnqvtg�?�k ��Os�\]�����*i�壓��:5�r$ Z����{;dMOܸ���Q����y"N��Ly��Ƨfy�ͤ��;gx���1��fv�>�f���GX���MNMr�*YT/8�"7UGk�8��L�����y~�4��K���^��		\й����ǒ�p�E�:�&}�cc,I�R@@<��zMg��T� wq��~x�awF`�7䳺��AS�U��XT�P�>��q�S���g��GT<��l�f��f��$H25��f�암dT֮� �9�=���(�[��p5��
Պ���٨��_�.؏��{i�����R�<k>����`��JJ_t�kH*�!Q��h;N���R6b7���3�g	ɑ{V�q\��TD���y�s���ʹ/cj��ۉG�Ve���p��X��yԋ2��0��|������5��g����Z�8��9�lt���4����ťڹs��� �y/�V��h[��k��X0�k�V�GhX�(�o������w�ʡڬag͗+������Iv�z<ي�&�4��;��5,T�h(�B���CI� W�(����i"�(!�bF^�y�� ���o�ɦC�`�!A�P�E��k��N^���*����d��OId�Bx��2��LN��4\i�*ʂ�UE�����-��Ih��Y�6:6�UK�~gMd�� O�*����9��j����7����ɢ���ӓ0�zƊ����=D����Cd�\�J����a�4$���̚1���;�d��&��tB�������4�� +nq���܆�D��M4�*%m��1S�ejU�?q�(�O�W��s�-�n.]�h���4t?�8�H�j4rO��P�Pv�S��{� !er.o�	rɶh8�_
��[�k��y���^�r�$������i\����K��,�'tV�* �2��_<Ie���}(Q
��>W��=�P��^�M�Sk��&�X��}���êK�t	����(� ��i���J-+��c�����K���]��]�`�)�mTJ �n~t�U�W�����VG��U!J�Vx���t�:9�.��cw�`��m۶ ��<�@~Ԃ�<��p�qr${���M�NR��B���8pM��5`���P�������j9�~�+t/WI�d���.��W1�z��E4p`Ye��\�UT��]K�����&b��
�+����S*��#fan��#Ϧρ?�H����U�X�]��F�PE�D����#�'�,�Q,"B��MM��������)�,{�A��]9���8���'� �� *��4	�/o���і�#у!��y�-VbAa'6j��6�MEՌ������8p�0�� ����<`��͓>[��;1=̘�Y����,pQvs��h�n�V����=�2�"�0�aŞ||{��SfǞ��nx�,�����fyn����+�W-��	�j`)Ć�'�yz��9-zp+JI�z43L�oX�{�=�t�o���K�+�4T'|��|�G�v������
d���QE�4�I���#�_����dBU⯱�i�3r���U���>fm6�d��M�xzo��A�ͪ$.!6�<^�[�4�W	�ZZXД���Cd#\����$L�~Xlkx�uM�*�<�:�=�Ծ���	B�Bkx�1��YԢ��H���򔺆��"/�,J���%s���G�G~�l�۶m�[���ì�h�v�FG���H�˰ú��*�Y�i����]kI��zI\���>k����8��C�x�JP\�4#W����|/v ���p�d1��+eI�03�j���G�v��yx�"��Ѧ��Ҁ֎9BO���;��˗�_v<zH^����M��J�t�2��� �\�Kb$�X�}K��i�P ��^^,J ���6\iQ��#��T���.�s��$�x�:6�7=�����x��gh�P,���f�(q�VH�ر��ٽ��u�13=�݂���n3c��5F����c�2ǐ�	��j@/�(X��B����t�q�JX�i�D	��=�~NY�k ���~l�Y�ψKk��%X�#�}�.�{�^�?����kW����͹����S'����<�d��>�e�&$�ѫ��,~z�p�"z!��f���_��B�����=����b�����XUx �L�E�D�<<��x�1ǰ9�� �@q`��	��F��m�aSV���]��+W�,�aװYӤ\<��"5��r��ʪ+�J�F�����J�+�O��L8U�Q�A-�[lR!�����9��@ω)Oҕ��Ρ�WO���Q�(�3#��kbk}p�|&w��>���5�U�&kyy�^#�䭇��-ٶ �-�$�7��^8_���y���$���ۂܴ�@a !�eV�5hhD.7�;�=�t�f|l��Û�4f��w�zr�.ɥBɖ1@$Ś��J�5	G�j��� _�e`&u�M��DC�z��N��lmP����Z=/�뀍�t��b�p*Z�h ���XV��۴��%���X��9�}vk��*���b���Mj2Y0��TZC����R�p��1�����T*������L�g��&�'��/��λ��("�ðxB=1�E�)�l���=��ȸ�����D�{�g&4��[�<�s�v�H�9e���^���) �b|���E	Io�0���6TԢ����g.��MS�Wy��T$��u#w��2䠊�b���d�
G8�^t�eO{�ۦ���#w�co���w����ČPX0-H�Ih����0t�)�&s���ՠj��&��f"߅�9)
a{�WD��^�j=�xK�y&�+c��^�>�R��UN&����؀���뙙]�̶�;���~'�\�����Ι�׮���yɾw����ŋܘLM�׫5�Րc�7�ࣣu�S!Ҭp�nB���bK2���v��岇}
O�EP&�o�;�����.-��y\!��d	ۃ�)t���
�V�\]Y�O�7r��Ce��o
�JU�T�sӅ޷���/�d������ׂ�B�U�k�Vlqo-H��R>����C���D.�E%�O���i�O?����H�Ғ�����mS���p*�[0�}�\�;X����P��ח��`l�yL�87E�>>۱�R�؟��fV�}�H'u���rd݈�k�iC+[|��}'�@=��ht̕+��|�27�W�]o�[���h�Mh�QAx�n��v˶-�{6μ���ʵksF�BoCӂ�0�$$����y�Ev=ߥ�	6�I��/x����ͼ�*����ڰsĥ�3=N~^�X�W�dף�$���*� W�*%�}w�;��-�����7� ��������~ꑀQF55xG`p���S��o����H1�U��w��j�W��IAH��*x�]7h���� �)*P����".�E8�5u�^�rB�,x�=���$�G"K˫.a& 0bx��`n۱�=z����̞��;ލ��`���1�\��S�G�dV8��7���C��j�s��O?p`W7)7�*u�Wc�B�h��C{Fk��ծ��*��H8��I���fh4/-�p�bH�۹o��޹�Ʉ?�5W/_!�y��'��?n�_��H��ԤY��������v,	��+ݨ��]OF�<g6���dD)n269N��� �JX^U6$�� ���i6�Y���j�˰��aǿن~v���%�j3��#���縘�;��_��j�tr�Q�"He$�gG=��Ag�NTJ=��7�~��_�l��HiHe��d�G�6��&��2��\%d��<���_v����X����ͪal���xo�&��)<g�gR�J���4W�l��N�J���NAAy����\C�ZW��ￅ�>��Ʈ/��¹���I,��Խ�5!?���5jb���(��Psm|y�u���ԣ(3�3=C��7�(���Ds�8>,^X�Z������@'���h��8����yYN)�n���%�)|ک�i��[+m��5��/@C����@9իW�2LH=��$/2a�U��Izq��]](7�`�7T� ?��4a���4�t,m����ش9v����cw��~�ы�m���I������x� ��{n��1����X=�&h�2+9���� g2�9P+U��Lg�z��,�j`A���j�i�Ԕ�n��*F�-��a% @F������ڶ�.����)�f�'F���ċ~ǝ���2���'��Ԍy�W̥K�͙'XQ%V
�`gt�@rbw�x��d�` �gQ�
k�B�3�+��}W.�B�=dIq#�f����6�0I%��*���(S�P'�,d5��5V-��f���7��@�2��P�Ֆ�1풢�~�6���i���S&b:�+l@�78vV�,q8�UoM�TJI��� HQ��ʟ���[䪷�e�f�p��qNXI/&�y8�Mh(3<w}λt��������u�l�߶xo�沚}��y�iGy�Q��._�d���"ߕ���լ�=��B��̸._Ùo��I��j.��fIJRU��Rτr��F���݁Ϲ��"�껌x;�ǫז�fo��`�n�L�-&��Z��� ț?�?̫QxO��H�+�ecv�6Zg�	Яv��"�MϩIx1%�b	����1����E,�+�m��'���`@���{�46���Z]��������|����s�=���m�(�:�@"*�)��N%��y���#6��H�U�����>n��*����5����x|�W2����4�g�*����L�pU��|vT�_7����ѳ�B"��Nr�Z7~�Â(/��O��(��T<ङ,���������_6�|�#�{�;a���g���0+(]���z�ǖg.��Z�y}�V��$s...��|��#L���N�k}�"[8k�3J�8A��<o�取و������Zn�D�cA{�#�Q_�=�Bq������y�WbD�u=�E�t�$��{�D��������Y�w���"K�,Y�\��B�z�Z:��4\ъ���/v��J'�����z�������j?��xo�����J�R�4�r�x����W��Hv��ur�\�E�ި�W��))��V.�B�r�T�� �^Vʞ�@6	3l�<�,��.����g�D�H�
�g�q� p,�=G�0�d� n:>H)Ԋ5���=I!)�t��o,K�0y2�Ã���ly�1FP/�����U	:=��̢��iLK���D'�_�@����x.�,r���	�� �c�d�����0�hqn!�"�c2`;�K�/���T�o����y�63�!�
��ݗ����C����K�u��jj�^g����bq"�2W%��$ʦgf8�1o�\0+�������-�|a��&��v����R����*9�MrQiIeG��m���o� `wfvF�������ȅgwbl�󒀻3�Zx��s�R�}�8�bд`�����Ơ�3#{�]<��t�-����.:�����x��ss</�#L��}߶{������])/�7&����1�y��mFm��I�!##3��f���� T_��|��es��9>����w�y��G��-�}�<��S��4�h�@A�P��2A�eJ����������X��ϴ_�p�Ĕ�> )6Y�h�ړGsR7/�;�ߊ�F�"9�.a�0��,.qn�~�o����A���w<~�E=�n�ݯêKk�{�b&�J�[&"j��tps���nU+�O)죗'煡J�$:��a��[^ILTh�z1sA3�{l|�\EJD
F��ot�!���x���R�&�a���D�"���Z�P������n�L�~�n�'r�#q���SM�n,�9EҢ�y���0"0�(��^$�(]���Dt:�$�?>.�q���6W��gNC�~�(���}��� a���j%�a�B��9���&�����\�rгY���l�ם=3��+���d�P����e]uj��lV�m� ��#Sܽ�����*��p�
�qy�w�-���P
�΁�-�Ô5��-p�v��H��e�P���
����e�T��î
r�uæ$,����͛^|��ع�����ogϞe�1�V{����Y�]K�aD w���M��0&�y��?�3X	��rf貟���Jvm�V�,X�ٍ{�Sf���#w����wA$
���쁃�j]�(�ONh*��jj��?�{l���ط�Օ���2ׯ\5ׯ^3��F`uiE�����3e_;'����H�@�&(h |��x��K�l j-�Z��V5�}�y�-�3�8W�����qp��[�J$B`��p��I��%�'�� $nC\��Hc�U�$K�cb�X�����G	�?���o?g�~�)��k�q�M�LY��h��R պ9�9z� ���
�-�����p���2�Wh���kv��{KK�%� ��V�[����hZN7�&��S�+�p��2�`P��\fN׃,� ��8.hh�V���TU�ȓ��Ujs�2YG�'���"�bJ�f�+�k�@�z�<e�W���]���ˣ�w���a��m��B-e0�6��[���X��`2|�㱣_o�F@C��i���L�(OWB�^����J�A0
n��oEqf԰C/r���9^p��,ox��ڠFh�V,�0Lfl3�1�K�뜃՛L���:n��Ev>'���	�k�&�q��D3<R v����p�c�/�rrŰ>������9s欹뮣��>���W�bΜ>�2���..ó�J�b�hm{�n�)�f�6��W�;^슇�(�U�#�+a�.�D��=F PX�>x��:l��s���y����0��v!=�kP�b��;�4��QI-�x-����
㕶i����նY�zݴ����kfuqA2��f`��A'(T9��G;�Y.u�R�Ќٿc,�=��O�XmĞK6=�h@�;>$<ē�$���h-/����U���Ƃ�+v�Xp[��_��m�w���f���fj�6� �TS��! �x��iUaC]C&�}?$w��h(#���4�� �ڵ׼�v��9q�{晧�i�}�I{���NV|&{��UzL�	�3�P(�6d�f�t�i�}B�F$�1
��s����&�ey�Vbċ�Q�8�v��'E�U����h�o�ߨ��4����}P��"/��k��<PM'ɼʴ=%%3&6��^s�-ؔ� ��U(���妛�|Üs{�Ѥ\�c�智��>�CE�L
��j��������Wr\�8��S���X�G�.J���q�.���NMM���CE�b�A8 d�'����bD6�>��S��zza�b����%I:tqb?K_U��2᨟'<�*^L`��&�|�e ��#4�^V^SA�3��HfYͬUln�1{�8�w{l�� �[���_��_Q�`vz&3����#���p��F^�Wu
�n���%m�A@����faa��������́�s�=�U'�lyzY�8��+^Ƿ,����3�nBQ�l:�2�zs*u�7fY^��4�c�ѣ������w�ˌMN1)�	����R؄�HvN7��
��+��A�j������k����+�����/��O(C�Rd�ՉF�
���QQq� w j�^��PH�8�$��w��m�����m0�k�'��bW9�ﴯ'��\��IC�L����	���\=w�����
S�ܻ�Lo��2�ԶY3ը��[ܵ]lCrlq����f��e�=��EN{�[���!�w�~s��Q�������O|�}N@cb�m��({3����[[G�HRj���<vC��b}��"������ݳw�Y^X䜦�}O�ߏ���u�M�jPMʃ'�&@�ˁ�]?b^MRq\�ܻ��w��:�$l���H��(}��I�i��L38�g��D-s������%���7���u��W]m����\����Y��K�f����oN�V�ѷ-�{�5BF�h��1#��.��9h� ������J�a�ܓ��"àX ���`3��`��]��͈O�A�G"�]	�B+����B�'�F?�9���j��O��&�x��c��D�!緒��y�@'��.4M�HJ�k�sQ�3�>4c�)FMu\��p,�;�qcU��2�/�?���O�C��Sf΂�^O
|�?eN�xÂ��vS3c��D��+���_l&��[ ��/X�L|ً4  jdd�ΟEr=�o'��ݴ|��6�=��y���\����Y\\0�j��J���Ք�/P"��l(�wj��!e]�X1�%�{��R���E^Y����؞��3��Q�x��6?����>ʀ-����Pd�Ȝ�T���V���R3Y�����KW���'O�k�.���s��Zd(� �X
�#��G�'�l�Y�ԡjBՎ�ſ�m��~�4�}�(7�1�@֬6n&�}6�	�Զ�ē��@x��nl ��$�u��-7�c��hM�΅����<]1�j����r�\_xݜ�齝ٹ��q�]fǮ]f��]�b�Ჽw��bzv�n�!l@�M�R�c�I�c�
n���>t��;|��9p�<�ͧ����Ҙp�P�4��Q�Dx�����.�S�l�P��0�X9�TB&?���Y�'=(n��{�g��H�V�r&�Ya;�תRZ����������J%Cr���`���5eE�A%O>���}EB%'�酭���oRo�Jk:0�)N}���	��uY*7P�n�(�T/��%�2A��L&�l,��#U�`��I���@[�Ġ��Z��S�W,��5������`�g�=>*<j�� R��A)A�6����#'M;�W��-��r��0�yP�sF�14�v������b��$d��w0߷�M>����}Ϸ���ϛ)>��nݶxo�[s}n�n [��E2���aZW�-�k����.|��_!q�w!G����Q�����p�5�x%�x1�ˎ�������4t��;��M��0	(����҂	�:3��s@]O���ۻIu�r+�x�z�B�������/s�f={M(r/�	�	���~��<��
	�ʎ��W��fvv�4,���s��|�y��������RUwI
��؉�0�s6�+"rR*x�B����q�7|BL�����zT4謶�]�{�:f�{�s���f�.Z�q)��m߂��T*��F�.��녦Y�r�\�x�,\�n�\3K��������[;b��n����	)�f���=��M��{���;��,�ݱk��ݱ�-��U)���Mx�<e�4d5�I�vS�Q�6X��~���4M;_�o��5v�1�����-8n.������"!�g�׼2o^Y��y����ܱ��:rȄ#frzҌ�ϭZ ض�3v�9
��0m���֫f$�H�E;�m:�q�n�f�ѻ�f������^zɴP���خ�\4T���r�C�)e�5�+U�^�Fz����+��IY�<�.쥀�(+��{�*QI+Yq�eC� �F�3����7�9!�`c����+%�:���
�+U�n[A�������X�X�\Oֱ�k���3��?�N��U�%��%��0.6" c���ƛ�Mjs\o|����	�i7�h֞�^�~}��w�G��j?ضxo���J�g�V`��#Baؽ��D߅��8^�8�̘#��7�bY����#ǫ\_���������/��Fd^�`W�qJ���L�r}�@orsFJ����1A8��ɒ\T� �^�1�-__y���H|{��1�?��9}�kx��5	��
�q�rņ�ɢ�_�n�I�^F�w��!�#���nA`��Ç3����^0;�oώMo
�.Uw3/�L�H��ɀ4ސ��fZ���jn=IΌ-����Ĥ9��;ͣ���ٻ� UP`��l2� ���]�ۥ�}��?�X�����}�Pl*�W�Y �4� ��h�1��;�,wQ̥c��5�G��N�]�X`=�{���6c<H���Ô]0�ݞ�#�P�|�[1�Ӑ�z�	�M+�(�K4��[�I�9��$��S),�� ����g?�c�����9xWO�1}$�<��T��Tj���'�����l*�Θ�|�[f�ͽo��9z�=G�R�=��@ ��/T ,�&p�R6�vΌ����������h��կ�W^9nZȍ�L�Ml�޻���OP�bq�g(-cѨ�?�Ͷ��U�m���.�q �Fb%���<�<)=��e�
�;�ܬ���9��ì�jxv,���g���QQ'���RS�!�������&I��~�wŉ������6�Z��Fzx��ϊl�\��d$��կF�݅�u�m�+�����F�Rl:�9l< x����\�(h����Gl?���5� ��Զ���`5~�3<�Lnq�Ȳ�����ᗢ1(V��C`�Q��a	R7� )���M���z���n�Û��4���Y�Q�����U!����f�^�TGS��x�Z�D�={v3���g�e�q��xw��\4�7qK�*	ϭ��Czz����ݳ�E��\���Vr!''���={��x\I��2X*	����樸Ж��O��c�T�ڻw�����̱�4w����4u����zp+��H��;v�Gv�}�z�9��q�^2����49>!�b��i�ZL؛�׿g���e�Z�^s}j�\mY�h�-�D��x�*�/n�{WK,l���["yU�rS�3	9����{�3�JjUQ^	ݦ��Ἵ�k�n����g��ŦӋ���K"�8r7��ՖY��fN�<i.�>k�)���ر����^0 s��"U������W_3����:z�l?��l߻ӬZ�ތ{f��`���Z��mV�9=�����͘���������O=m�y�is��ݼ�M � ����w�Q�x���s���4e!���-lRI3���!2|�",$UZ�[����C	_�� �k⪖.g�rԷ�U�$>QIm zc�5����&PCQ��F��� %����t��I�s��5�}���q�+R�X�H9E��BF�,h�Cgfzƿ>w���g������ཅ���+u����~���( ��I�!��«�����S�"@3gȱX+�h���	�wVE��>��F������:������^���a( P���n��T͒�%��C�ǆ��B�B�S�&QQ���T���8,���X.��R�R��G���߲`)��ڦ��!c�>y�I�ʚ�LH�^��2x�r�o��J��m۶��Ǐ�v��}[�@IQ��qWn��.�����+{�a��;V��>��	R� �Nexf�s���̞��8& I�v�✃������,��T� �T�+ln��x�HhcQ�+�p=��h(E*({�"�X�ٱ���2��O�w��3bAw|�4$��Q�,m�y܎�x��:b�s��汿��9��	�4;�������q��I^\\6���TA�}�!� ��I���^n��h�.^7����Fmzm_��=I[��p:�- o�w���v�=z:�:���n"7:�8�xj����x�x��$����	@�=W�����̓��G�X^x�u�3�_�h�-� ڥ�>c�F�g}�vꜹp悩NM�;����{��]Ӧ���h�v[�X	�=���Ȩ����=�"�_8df��͑#G̗�x̜8��0]7v\��lR�8��t��L��������R�G� 1V	$)����}ͰGCR�m���[!�� ���u���Mm�$D�緘��MA[�IPN�����a[I�c{4g7�Rr��pv\�염�����2������Ue�0/��g%�I`Ң&z�ݤ����U����'U �2S�}W	�
�l���͉r��3�����\�|��5�!�������޻v�}F��jmP�}��E�͌�V#e�A�'��Z.^���A��\/�-��Ҷ �-�Z��X�՚U-JY����!9���`k����Y�b��U�K�yV�li�x;��FAF�P��U+���W�y�o6+�X>N��7�N���"�QR���{�N�P26k��3��
������>����^�S�ٶYy��iW"��4��=����C���>4��1 (���HnØ�}�n&��:.^�H!x.va�f3��m`'��$�~��a��-3a��=�����2G��c��J$Ca����h����Q��Gr���s�}�|�����K��ĎqÇ��v�NŸ�+��8�k�ٵg�ٹo�iLL	\v��a�����7�P,f��a .�N�}��$ͮ �#�ƃW6����@l��Ķ�+�Cѣ�{I�%k��J���}��.5�,��\��v����������c&�����ݤ?���	��ks�kǵI�7xϣ����ŧ�y�\z�y�=������m3fn�h�<6��7��40Kv<��&����y������0r�����y��o��g�$�u&x#қʬ,_վm�@7���4@� -HJ�$�f(͎���Y힝�=�cg��h��hVf8:�'EI�H� �=ڡ�]y�>3����"#��� �D�U�PU]�/^������}�#`����6���eS�D�]��8��n2�И֦��،* �,¯�t F]���ڭ]!�ׄi��.�}�����R��2���Z�ָ.�!�3�춙/M�������(�k5�o6�,��/D�s�6�e%�<�~[��҄�θ0y�<=]ik0/\{$A���1"�y����ŀw9�{��e�{��b�x���xL���2�Kԭ*HeZ o�%u�&����QQ0T���kc	I0�X
 ��+ޯ8�пl�W�`���Y����v �f
��� Y@���#/G�آ�E&������,��R����)��e�^,H7pO�'O����p�,K3�����)��w; ��@d 5�%x����|&|M�\���F�dӢ��; �!=6v
ڔZ�?"NY�|����Hͻ
���Q�im�>��. ['�]�IB��GV�U۶�]w�C`7��0G�����Afʆ`>T6�\@DQ�R��/lM;A��$��a�G)�&�1�R����V�W���P�5��Y�D�d�`!ܕe �#���TW��G�oMΡЕ�Q/��r��RA���~��ZH���q�<��G��7V�rh�ku�9�����/�����@���'�)G�]F����9r����"-��?$��i$md_˔�2x��6-z�?�+����]���GD��k��e�Er]����<s���o�[1�r}�_~�?y�N���A�M����\!#j�o����:hꇥ�K�@��,�H	�ZTK6��Y'�5���nD��; ������tW��Ţ� ɀ"���9q���M�.�9��)R8ii��ߍt���V�bz����&;u�+��9���0m��<[��N?����1rB���de�@��Eq�N�:e�]�v�^fm�^RM2!�NLL؅^e+�[�R�*F3�Ƴ=����=;i�a1�9���t�Z��i��ϒ������ۋ�̹uN��Y�~�ֲY]<�#E�f�˚-�6���譱ֵ(qu�<�� �Ȑ����[�Q��~r�����V����� ;ԚrM+V����7�������Y���aC(��癙�@�N26�IV�� ��3���LC�c�������t��ӭ��!���sӲ�)��3Ў&���T���e�y��}���7�9���l,!�k�x)�i�5W����~���!�;� ;� �ǨEM�1Qz���呈8���`�`W^ʋ[�i�S�s�a�M �dnG�N�uT� �SZ��xB���x �8�
H��_�c��fGE���xj{8�|v��y���
�l�HG������S�A�	G�T�$�ű7���#Ǩg������a��m��^��TY��Xt�<F"���������P��~�^z�E�	 ]d�2��Qc���Dh@@7�i�k�Z4���M-�E�,�HsI1[��u3�?݋]��[Dg����Ɓ�N� ��� ������΁1l�t�����eQ}��4c��Ʈ����i��AM�~KE%P�	*
H�="%���͙v�Εo֔������{�R����Xj}]Ƽ�S[��P��ω'�*r���cGGD����ߑQ�TfP�q6����L������:�����n�`YJbJ�Mˋ�)"S�Yg�(#S�/T�WU���ō�0YT�Ǣ�D(́>#��jSf�����t��oD��� `4���4m#<�,���zqn�����<+�^�rM�zI
��W��ScTnT�<!��5\)�j�cqM��@�ee����Z9lڴ����lg�/�@�9��S�݁�6\ C��07t���t��~2���j�/�hhd�~睴f�Z����e>������r�������5�{k�-j�W���^ڊ�xT�����^�h�M�#�ҙ�����M[��{�U�׊�.��QP,���uŸ�Y<^�uf6�9:��a���kt��a�3hK��[ՠ��.�dˆ֮�+�l&+g��S�;����D�"�F�_��y�r:�uq'X��o���5j��0xV[$�� c!�{I��m��ʃ��lQwh��D��G� �8?�&z��q_�m��.~��{���=
 ��5M)(B�h���b��4�� M<N��N����r�UwE/�29KE`S�ǩg�m޾�F֮�yˡ�fU������C��f`��K�E���n�6�v����48�Oc�ǩ`H����0����RF��!����X�?Qxf��&ȆE�/�~ �h�Mz;���k�����#s����l��+���ɴXj�>��gq��1�7l���Dx���s��IQ��3�M��:`�l*�����g�����S�̟U
l��b��1S��$���q���-6%A��	��G�k�_��E��z�3-��)K�H��{�� �����䞛9��3�KQ���(�GN(,ZZ�I�P�,��@%B�\'֯Z�B�zB2�F'Z�^�p�wЃj�eR	��W-A�&n������ז��,�[�(D�q*+46vZ���PZY�UE��]M�02_F
�h�!��Jrڷ�x)�0S�k2[����f�lY���]L��޺�lP��ؙ:�?��t���"P/l%�.�__��;�kS�iC�ʆT���*���h�����6P5�QZ�z5=x���{�>e,��� �1��9G� ���t����*�V�N;��:7h��9�/xzv��rݔ�+V�g��E)H�@��;#�NK�����'�� m�3��{��E���$�rn����m�zm��J�wS�4������}n"�WW�k]f�h���g�Tx,i����&`	�*���y\m)K`��x[a~��T������dN}�o�)2��� ��5��l���h˕W	w����tt�~��U�1�����у�h�݃�����;��1�0����&1lP���ܼ�h�4g��h����/�6���~�[ߤ1�ɮ��p�MMS��]�����|���%�'˧�2�"YE�eB&϶�xU���~q���x�;��9π:��>��3��>2}`v�>Lk��/�_g���d�V�rjl�r�ؖҌ7�b&���uq)y��b��a��%Шv-\�}�X��M)�8��_F��[[��Vc�[����\�r�T&L4�����`�� �ᬨ��U��mk��!��ɳ�aL�n"�̟�����F�J�e�/�z���F/<���]U�K�=M�p��y���Z�����g&fh��y!QN�l�"@���q�#���+�����h{T���R��=���
�xu��2Z�ԩ���Ԧ�������Sv�:ۄ� ��_�`�P�;H��{�vd)�[#�C��A?��$sAFJ�_"�l���-VjB_��#��> 277+�I��z��Z��Ki�\ɥ��3z��ש>_�|2�`Уj�BVâ�:������շ�@n.E���8%����]B������:M�Sba�w@t�����Īp�Bק�{�a������D���y�6� J��巫t�wy�e�V�_^����sr�s=�����6[�T����B}�Wњ��� �٭����s|/�T�+ҋO<E��K���ߡ5Ct��1J�ԟ��ɩ)�൸��9b�A-���u������_҉c�$p��F��u_�������,�6Jޯ�ur��ʸ*�/܌���z���VW�iT�!���'e�K�IQ���R�@p�T�m������ΖQ�u7S�f� ;[�*Eg�FK��n�泄�b�b���@z���x�L:�aL��b����}����Z�j�����hˀ�jx�y�H�c�e�D�����n'�B>�-n�dj=K�;s�m��-td��t~������)�k~�[ ԍ܎�Fe:aơI���MK�BcP�	�������&PlQb�:z�����ZS��ί!�nXP��v�}{�R��/�v�hXlatn!�GDo�CM��!��4�Ʋ�G�c6E^�ne&���mw�I;���X��
�T��#������T���z�A?���ș,�ßcÞ9������b�`��{v���5Խr��l�NW����n2 �D�+0��U�s�A�I�(�K}ϔ�W[��S/|à���.��j̭Ƨ����dpU��4�m�� ��Y]\+��0Ą3�ϰ��E���`E���`W��m�/��*����������òuf���EC����}���W����hݖ+��ic�ۗLK@gs@S� EXp�<��������}�������������cL�|�A9_��[:�n�&��.E�R�X@�H2F�i-�v1��}�]4�Pk�\`�����K����-lnn��H�5sdˌ�%	��]gy[�6�Ʉ�$4�3���/�i�תi�Z�;��^ Û�`�Y6�����ݼ��%�4������-���>��@�`dH:�k�P�����͟Y��d��ЎX
	le�kIvEe�$"���T���L=	`r�OJ�[� ���]!Lb8��`��WX�\�FÀ^K�{²A�/�B�V��L���=��v�x�����\a��r˵�������a�g�սP�j5�yp!����W\��&''�= �bs�*�dc� T�p��9�hK"�
s�a}�OS��
ǁʁqX[�z����{�����Y)2�y�N���y�K
���S��N.2� �F��i�?EZg�e�Vk1�'�^p�a�P���>� �}��D}�T��
�x����PW7_x���1�(�N�3?}�掞d��S"��d!GE~&��G�l�kn����XCN��˥�f��\�k�#$�
�qb�m�Կliڪ �Qc)B�ͮ{q0��V�C�핝����8�{� ֨kؚ"`k.�Y��%�����Q�6E@��{-�lָm���M����\�J]Q����vڲm�{�mݽ_\�2�$�kUZ70$���������N����L6O��"E}5�<ˑ�7-Z�.ո�w��!�v_������x�0ehR��q�I�=:s���&�!�ƺk�
c�� ��=stf�B@��@�E4����y��'O�Kg��(���B����q��3Z�q�yu��)�TWY幁��3�fF�o$Y������"=C%�Z6�W9��2׉��)��4�1����)��PiYL���4����&e�hL�ё�q[�V�W�b؈��4|n
�Z�\��� ��%e�1�dW�S)�e���O:����x,d���:L��7�-�K���hU*U��  BL*�A��t�5���$��T��b��V����;�������*����m4�39g6L�����դp�'����R�-�8a�@^_ƙ cI+g�MU�7Ht��cLI|���P�V}p��~k!4VԘ�{�42<L=��dy�m��.���߱�?&��eA�XG�^Mq1Y(#a���*��Hă,��B��w��g���c>Lw�s/�iC�lR2�8��6��/�%�\���}�^y�9�5}�Jx�|��F���z�]��Pf�|ʯr��ͦ(]��E�6��Ѹ�&X�q�,����S)zY$�, хH
�B}��v��b@� v���^���j���o���0��l(�~�Ia�4;5ί�Q���n��Nںez{�6�����N��}��׏�?�m��::57%
�LR�W�ר��8`IIP�q��.�p��}��}41=M]��Y5�k��|� �
�[�1hJ1"A��3���T���MC�2?�r���s��e ���P禒�%(P�Φ֢h��p���*=G�ZҢ(�g���k��u�[x<�/�^����X1u* ��'��:��%'i�]Vm�^Z͒-o�hGGGy�Vَ��)&���U�9���L���_������H� �ҙ^��tp���IY�XLɺ8‣�l���_d�ZYe[�k*�h�R���rF��%����jCd15�W�	�$�����g�ey�ί�Xdl��vW�^-�Ļ�|�*��=JX=*`��[n��;w�{�G��C���k-��r�J��� �M	 ��U��A?/Ğ�@�u,Ke�햁����$�Jp�P����m�z��e�C�l�=}��`�19G��.���hϮ����Sw�g��-�R��y�^1H7츙Vl�@��MGy�1ȅZ�VfpV�E��z�8�x��m1���f $���U�.;��Rsz�̫!�����~]P�%,�B�^�|�y���`6x���-N���px�f�<��TYFK5����N�$��4�����z��x�w3��`�Bc�R���m��:ɦ���Ej���OS�/t����=�ēt����޻����92�EFf�+����&�
���W,���y� ��:ߥ7^{]����<8�1:��/���#��w8阌��gV �h�"(����NP�dcb��6� M����~X�*��j �-�>�~w�����_(U�3�ǒ��"H��s����]�Ͻ�2�h&!�E��X�+c���}��"Z?��<^�#���mj�Fd�+���/v8*�_,sx/��x/���`%�o�>�)�T�QLȆ �腢Ӆ�oq�Z���j�x9f��U��� ]D� ;K�݇ut#3��L�Lh!��Ų`�/3����H�w��� �	�S���O�q ]�e�5n1g"��^�1�ndUGF�W^����v-ُ�������:02,fC�� ��� ��ȑ�K��d���DS(P�$���ώ�T���D�-Wӊ[C_��P*>��Gh��*�!��J�I����85G��C�F��������{R���P��f�稙�Ѻ��҆k������r)�jTD�ϔ��q�Aف�/ΧX��9�c�eq&�=��m-i~�Z���m�{;?�s�����l��V�Y�9T������R���J����n��	Kk)5K������{P�}+]�|T��c��Q:N�G��������{ϾB�zC�6��0�6h��):�C�ﺝ�ɸp���TjU�)�3�N���o3��i�f��/����7_U8ݝ�=s粽dx�ֶ���F�~=��X]G�8�@�cQ�N�{`)ɬ���a?*�-���a	D���os찎x��i�y8���S� ׈��8���LS"J��	�.`�o�u��>X�"r�h���b�(% y� 	�~����o��G�T_n�-�K�)aOfL�� ��2495N���T����"U�F�4��*�0[& #�d@Wv����ηc���!-ٴ��qJD�T���J=K�����X(S���d�xQڻw�L�OPWwVx���=�(��[w������JIT:36���:()x���#�ʊ4��������Յ�zm]�k�sן���/��9<�a�!HpV+5j򹪬�'\ئ�HQr�˪���Hp� `�bx��?@�܏�DJ�݊��EwUo뙆�������{��T���U��"�cL��Y�Q ��D��ȱ�T����g<ߗ�r�+���5}�� V�����̮d0�6� ��'	��ʜ9���Q�j��t	ؽ���/�P��gS_[��įr@M���^�����o�$����34]�m��*�r��Իj���:M7��g�� �`�c=X�J-��|����`�����ؒ<���.����څ�g�W�S�C��ӢP+pi��Q�
�X��"�l�8W���
��*9���%�,DI���D%{兀�b7�m|M[���]�j����9��V�D�9*�<�Ў���׿M���O�.J�XX�i�D�o�G�����/��N����A��s���=����y�+����O>���<��ц�������>9�Z�H�TV4�Uq����ƿ��g5lG����J=���pk}U� ;Z�gƸ�+u�=���9Q���I�~qu#�ۗ�N4�9������H������T��tԧff��(6>! l�T�Q`�̳�����c"���{}��0/��m��и�Q��G�t�X,���}��E�V�rƬq������H-�����g8���c���usl��u}zJ�	��tF�y5�?c��,"�S&ӥ�������v��/�J�����s.�?�|Z���v��cD�������޷q#��z�d�w���0��L�r�Pm�^B���TD��H$���P��a�V\��G4]l��?�d\Ͷ_�������0<&2 �r����<i✥��[2-L$���zPHa8]�}�Y����Y����Y-��A�+���j�.d2�W�-�Y��\��}��{���'�mbnB�YVp[�(3����Z�?��C���2D�fC�����+i�T�J�Nu^�����y,�<ٗ�%Yd|����$�	'��b��5����Q; U��No��2�_����`��@���jخ������u=C4�� }�?�?��w�6�YO�������o��Wm�to7� �&9q^`}�I���W$���2����#|/��W��
g�:i#�9��%|w.@~��
�����7x����<��ý�\��l2`�R����c�w�W����)S�6�O���,5�Q��_�-��ɇ(5�+���(0��h��5����b�r�=��N��c�h��o�ڑ4�A(��1����)es���W<�E55�ٺ� �����V�٢����.��0>=���٧�&]2Κ�kv��m���l�Bk׬�>2��g�;��g@ �����T=�������V����Ai�۝����h��F��y4�v]8������e�{�5���Y�i�XOmG�������v6���^���0(�p�Ն�r3E�t&Z�6/f�(��$ q%&:C#NH�|,����da�>��L�9R\u�B�*k�ɂ'�et5��q� �]����|�E^�`� [d��>-��=�f��Z$-�MES۶�L��P�֯_O=�UQ�@�^mH� ¸�)�ݲ�m��������/�+]��:�*���Q��Y�ߨ��Kwe�G���b�݀��p
�\/�SO$I9�����*���B�X��N����>J�)�cj�5[��wP4���f��kuDg��aۓm�dz�#0t0YV�X4�v��3V�^&�У���2"Y����dLI �tt�񃶯G�٬j�Iw�A����r��Ȝq��je�(=�����<��PM�P�:<6c��e�y��E���#�)���O�������t��q�c|& �+N P�x�uF7�x�p r-O�b��s�1��+�&a���,�jS��@;�\ �|�h�Y����	x-��v��%��(�D��ł\����3�gjH ��m���wCq�T�����:��7��s�%��Oh����S��j�k�}��y0V*���w�^��vٴe�{	5L6 "+�n�!@&
�EU���@Eڴ'�$��Vv��޳1et[�	5g�����q�v�٦G������|�e�r����X"��!���=[3��L�D����v���4�ռ^d�����~��X<O��D��mI��_�7-%���b���.��-AG�˽��q ���N�h~f��Ţ�~`q�l-6u��3�2�1����B/���Ɩ��@|<��Ć[ωt���>�q������*�p�j�6W��D��|�G��Mo>�<1Z��,�)��E�I���:��3459FP��$~kPp�MsܲU�.��._�!<* �K���&��.>��4v�Ɇ���F=��.yB�:_�mJ�J�z�Y:Y���7^G�OO=�8U�d�}�y�L�H���C���(9P�gɊ�b��@�(���t�(O �_��/�7��t�ĨHR��_Q/ȴ�p�/�#Ԓ�RY^�۳�]������ò�(���E/��+Ь�9��@��/�h|���Y���
��%)pNn����K�u-��U�1Qx5��2�w�>���%Q��9�x�_�x/��x/�p�(�7j<�e��g}EIL��|���,��"��,� h,6�MEu�w��C�r1MEL�����~�p@�QiK�]�*Wx���QK;'n�%U��	e\ZMesU�dE� s� ���:팍҄�iiױ���k�X�n�4
�u�E�5=]P�P�7"�(F&{phP~����mY,Z(�"j�nAYO�jR��I����' .�A��=��}[�R�"`s۶�t����'��ɸ�p�P���A��Y�8 ��RT����2�h5�h��?,=��1
�D�NIT��y�~������=��$��"�\�t4E+�z��_�+O>M�O�H�z�zhb~�V�[O�=p?%{���8��&�zs����ͭ:�'q~/4y�j_2465��jޭ�rٳZ}�J��wd�0N-��/n~}Aࡣd���������m+���"�Xz�;��1�n��(UI��ʰ��hC��U���h���ֿ��\��4?1��~�o\Ew?�(���_�ܑ���c�(V(�N�sл�Pn�0Y�T��6�z��'(�0h�珞<NWl�L���g�����$5��S�K�ez�̥�쮯4�=�8���B$�Oɳ�g	�\\]��ۺ��W��؝��<9z\�2�H;"gjge���讓�����:~���>ʦҁt��2�#��������y�F�B�����l�q�2u�mJbR9M�z��-�&������lY�����D9Aƹ�	n��a�bd��df�/�߶ޝ0j��Z�2R��/�V<�v$�q�J��m�A���.?x.���Ж�%�\�Y�j�$��EjEghUj�O��\�35���8���S�H[��gv
g��w��Ri�V��� �t:����4�X��XP���g�y��ɾ��"��ZT_��������D���B_��qdv�󙎥�3������6��c@&&�2>@��ⷚ[M_`�k�����.�
�s�T��\� ���Qދ
�}��(Qv���&�D�?J;n�����'i�V��F��#�4:z���X�i���d����:7_D�ݧ�u(��]
8���'����.�YA��g���qe$���-��k5�w6��x�8�:�OBW�fR4���O�i�>O�����O����G��{�2:�]�4Y)R���?�!}�w�@��<OJ��j4]�q��yb����>gQ��5i��;賏}���?�%ug�d>� �1YX��d3�,ȳ��S���y��Ο��򙤟Q��e��@�E�F{��͒�7|��EE�"-Ԩ����õf^2�;��]�:�9�j�Yb�8��N �CA�m��9\�%@�Z먹��$2fV@�Jdl\���Ж�%��� �5����+3Tao�H�\�҅n�����baB�����!3�8�Zr��Z.dk�.�B688(�����vM��^�؞�5�]�@D�
�k<��j+�՜o�2t��믧����2 k�Lt=kH�Üh���	��D<��Bpt�Dk��Y�5E��k�-_U7G����ȧ?%�;H�I1f��`�K\�r�#�:}�=z鉟S��Ҋ��҂��Ц�����>ES�U�6���=B=�}Ba�>��-Y!dƚ�6��@QheLN�3CNd�X�5�1�i�й�z8�V���d�ｐ�s>�|��yu��e� ��~�� �j��nr~����(��i��t{+�nV���<J�l�#�<B4=K.�c��r� =�OO�#��EР� 0OMOP.�MIRc�ā��������k/�NSc�T�����*[��A�x����:����	
��Dte�� �D��M1�
�!>��������R���c��/����Y�qU������Z����պ��ے�gx;A��ɰ��,���7vϥ��}�[`T�����^������d�S�����b�����������e�{��e�{	6�@�H�j,F5��g�n;#�N�pvһ s7���ڸ�8q��C�z���s:ۖ�u���dj���{bZ�Y�3��2����)�+|c���vE�ɥd��֬�@{�A� 0ب��X�����Q1�Ks(ҁ��d�$C�Π�H`1��P�hQ(���g��s]�r\l��2����8��h���3�}��<L����\�Vl�H���4�`wگ__��{�_c ������B�		�[(\�愥����w��OVP���̮lu�������hz��QDh��p'pr�t�.nV0�:y��+�쁭�������Ȩ��LS:��D&E��\�JC���U���]����:�� %QJq�;}�4�
Yz�k_�O��ߦ�')���@6O3�
�ytY���"�4��6��?�ɿ���O�w�ǽ��ll����-�p��6Dg�7�,��x���*���#���$�խ�&�Bd{;��sQ�x�g�����DD/�|g=��toM��l�ӆ����`��Tv\O	k �^�9?Z�譕�j[|�Yߪi+fC��8qܘ_���.r[��PC��蕴U���ńSW�V�뵶�����6V�&�=���q�R�n,�}7��F��Ӽ9�u�,�.Ђ��iR��U4xX(��X�v�a��5M�#1m@��l<����|X�A�Ve�/����0���>��~�T�j<E�hB�n#х�dB*��^��x�B%5
��pV{�'D�Be�d��l�R�0���f v�>�~�d��N@V\Ll;9I�+V�y;t���P����ҋ�¢����;�F�_��0߇)��7PjM��2����܆�����1�K��G$A)��Ź�g|�=�[�%}��7(�4n��� ��i�����uz��'��\�%��R#��q�6�r�x<Mԫ�0-�� ��0��d��1��M����SkR�?�)~��q-�Vn�)�J������V�ązT�k�T��.�1v �%\o���^*�[�Q������g��M��
OMLR*�ܥ-T�L��|!�ЕnU�;����,�,���ldk��m��Q�*����v�j��XH��x�(c��[<�����L��4?^��(!��c7��1x�^$(q���X�?z�v���z)ʯI68(�-��]z�O˼Q�aWtWT<�eGx�$��`���?�#������
=�45>#�*h�� ��ԅ/���e�pÁ�O���69�������H�܌n7�v6��y�<�@K
7�n����~� ���=��3ׅ1�3HzBE®	vd��Ŷ�P��e>��`�}�0w"k��8G�y�泸���`M���w���v\����R
՗�5�|&uL�s0
q���
^�k:�Z'���C/:����e�^E��$d�M�s]?��;�״�#6s1�������<�[Ų���ۥۖ�%�<M��d�P�a��Lv��3��<-�\vNX^Ǆ9KTn&AOo�/�!�kap��+�e�>Cկ�]�$�-� j�-S|Ě� ���N�̈́JE�TU��B{���F���=3��<)��H���/"�V�Ud1O�4�ӆMW�]w�+��D*p��I��z����Ff���,�z��(��1��ˋr	�������v�G�l���^�}d ڝʑ[�Q�Ͽ�������?�9����~��W^Ao���(�W��T"�顙�i�Q)�����M�Qۨ�|L�M���W2Y�$��ݕ�,u�A[����g��������@/Y(޳l)j�����j��9��5Rm�(��+s��_{�{r��U�Ł�]�S�b>�2��$	v������R�7\H�9vEnPK"p��G==�$�Jﻩ�T��l@?�����c�Z*��#�I�U��}:1>M����o}��wh$W�����[73h��ǿ�m����4�\&)��@f>p@�pp�u�V�w�����O+W�e�"� ��U*5Qw(=o����r�֮���)Lqz[F5f�	}�˶7����j��2�w�\����B�����^"XE����T)[�*����]�s�&���6����������q�~�:y�-ٖ�%�L���uS$i{_�,f� �s�\�Qm�"?��8L�� ��F���`{�l���[�DA5��Zi2-Ov���7w/�ˑ#���]�� �'\�PAZx�9�]h������F����bǷ�����ЃJ���7ޠ���������^����딂:[0�@?@�*�!M
�|�6e�l�H�8����(�\��J#��Ў�g`ЃH�y'e���g�[<5AO���/�E'(+;  ��IDAT�Pt͍����S)�REw��GT1��pi���"�5�ݽ���U�&������'�.�;_���P� �r_t������;o�c��/~�,�Q;�Z*Q�vWƂe�\��$��j��sT����|�\���z���M�9}g7�߰������p�jT��� �*ܱ��i�-z�^���rKPbj���^�D�j;�Z.H��HG�󝙜���>��A���d:CP?���l"C���U�鮏?@}�=��?���#��Y��|�~��@�}�|�}m��p�k`U���x�}��/w=K�z�y���  &��P�k�gn1�pH�+"|�P�@�Nh��3�� ȅ%xF����q�5���p��07T�w�n�PE��H>����,�u��Ԕ���f+�҅?7ޯ��"�~q�2��k�I��i�e�{y�e�{�5U����?��lA�Fs��B���oI�\Nl�rW��yr��t�%��h�d���b�.t�����h!xQ^����aS��C{�,Z�w�J��k���Z)/�����'[�"�f�#�����ʕ+��{�={���s^O�  2�(\�"*��JU(��uu�G��[��d���D�'�d�r�'��'?N##��8ܞdgN�Q���T���[�^�����9Q�819N����~%��8�2H����d%��*�1����s/����T�e��N��R�mR6����<9uOh��:�x{?%$bI�/���ݻf��RE_C\����a{K�Y�H��g��s�S�63˿s�To2���������M?N����x_(7�R��5k�G�}2-\_�R�·|���XY�Z���L	��EM�K���p�T!\a[]ŧ��`[\t|~���ᱏ��m���s U��l\E7�{͍M��o�}�+�
�ݗ_�t6G7�st�Ds�z~�!?'aSe [�pP3C���J'N��C�ާ��7��#�|ry�Cֿ+�hWS%+���+(�^c:`� o�紵t��^�� uP�@8�T(���4��Vw����ZL?�L�wib�7���@(]�v��}�����F����~b��bi�S��.��x/��ɴ3V,�J[��e^\�$��'��bf��n�^�EV���x07�Un���3��'~W���dk:�Myc��(����\��/Ö���*����T�vپt�-S!��e�M��O&��r�,��?�Z��ز�Nr�vi�����F��m�P뮒3�n�:��*7��yW������� {��B���K�����@[��#��B�6@X`��n�3��b
 �D:�c�Dw�}w�[ˤR4~z�z{{���4:zB̓�G5\���>}�����q��_��i(�W��ei��$�#	���z��h��M�b�Q�{��d$S�#+ɟ�J���_�u�#t��Q�8޸�F��DU����
%���R+K@�ӝ�!gf�^�9:��n���(���E����ք�����Ԍ����ij0��2���V��c�bT�)Qib�zW���WW��F��A(�< cK�EW�q���4s�4=����4�]�5��ȝ�Е}���SO���/�"Y���0�r�f �2�r�(�,������c��sAoUޟ[%�ݱ440��9|J�x��+bh33;K��s4À~nnVKb�0�d!ł���p?�d��c���� �y�R�U��U�Ѿ}�ӕ+�/}��W+���K�f��<.�z�]/� ���;��83��9ѕ�S㔌fy�)��H ��g���?������T�*�8�� �Ȁ
�U
�|d����|���V]Q�xtp���X��j��&��P+��qUUx��O�s%�S��Os������Rk-��V��, Ö����*|DV�U�-��X��6;T*@պ�Z�\�i��є�����&6�-��b���M�8�x_d	t��Bh��1e�xL�"s{(45��b�h��,;킕[��nhg:����)�����D%�+c.<5�sw<��s ��s|֖ۥߖ�%��RX��a�G��%�MkQZ���c���s
|�	�5v~�}�;;^�a��b��W�*�6������9��{����iPB8v����B��Ƙ8�]����A
*`B`;�F�ՇD��3ϖ�)�|�?�iQ,�f5�|��t��!'�������|ժU4=1E�rEx��˝����l-�EG
�ܠ��4�﫪 o@��v__  ��o�����F����t<�!_�"��|2C��:@���G�<[ɸX����OR3��:��x���8Jr��?~���|�mJ֑V�Sůӵo��5+��� K% �4W�I����[uj���%�	J�0�I�,�:�
�u�.1Lm��E]��=�?�G���`�'��`a��ڽ���>�������A����������N#�+�����c��ǌ�z�rj�0H��A�VK�i�<^��;o�A����:yZ�p�&8�8�$SA���a��O|\vDE`n^�<F� 7ƀ9߅"�u��$0�D�����R�o4�� ��I@�7��W�{��W��~�%�a ޠ�tV�C >����f�5��ӟ�,}��K��>��+|]&n�����C�稫�n�.�%0o6[2l�	Л�����+؋�4_�{��*[�SP�����/������ԽV	C35���LM�	�E+3�E���hˀ�k�d�}�����\�x�m���>e���k��ᢀ��Aq��Y��-x�;�*�P�ťK�1�V�6$#��;@'���u�^�T��I�wgU�ݖ�EV�	ܓ/S������Z�F��|�8�͎MP��&�hp'&&$���]� �ծjBqp��������ۼᾎ���( �c\��޾M@gM�ݞpok�@=�����О7ޢ��I����)�_�/�Η�ϧ�ʤ�O�T㰮8?G���#	�yQz��7hߋ�Q���H� ��LQ�ֵ4�i�G���K2���U�[��͔��С��H�����&�	�_Ҡ=�+d���p�2�^II�� ��^}��T�:N�=���uq[�z-m�r]��
��8p�:�>��hKo��	�U�����fw�8�>���Iz睷�_�@��.�8qBŁ�ڸ�
Z�ne�)������|��������t��I������뿤��qڹ�^z����y�.@j�XF�T�$E(	D9��Ӎ��^��#��`��P��}�X����'���=�q��8I&�Tr�.Tt��P&�E���裏�k���`���W�Z�:�^�-���v�Un�������y���3Ƌy�A���饙��7�&�.�c@�s���49=�����I*\Mqq����`�d����j�`㾂�х��G>b�r�pm�^bM�(:A�7��|���~�dyC���Em^XP�tq���d��7k^��l��~�����@L�-t�}w6j���<�Fjg?�:�+Ey
���ߢ��UY�V`�<)�*�ʪG"?�0��d�O��	�2%M�c�1���Z"���v vv��L��rY2�F�M�o���w�r�4�� Pgp���{ｏz����2�:�=2���
��Ȟ��kϿD��/[T�G�����=J�n�20��U�}jlt���(W)� b����{�Kѓ�V�)Ue�w��M�7�O�c��#R�6S*R_:� ���ъ���M��|��gRyJ'R��"��a�^��c|j�Չ���8�$�"1�/��{ED��TH����Ok�M\s==��'izn�~��+t�-7K��l�B'�st��(�^IVO�? E�����9���������E�v�Ww=G)����Iw�u�8@��+� ���ƽ�0�ڻ�]z���k�7���}�/~����M�z��A�\�@0��P��
�ea�J����Ͽ�=�7�oUy,���y��z��>��B��yĒ	9���	�6'y|��_�?��?C�n�@�Y1<$�P�٠35�]-ūR��Jv�LN�xE61����
��"�ehM1�j����/l�.�mjs$B0�urx�h.���IS���h&� 2�g2/�&�u�
����2ང����(��Ji2��������TF��ZZ7Kج�,r<Rr�P�Sp<ɋJ �$+��B2�dc�6@$ A�v9Bf����'�xZ���L��*��A&���k9��oQ�e,)���R�V�b(H��!��i�E�Z�� �9_s���8���\#
�@���ڌ�X�����"��q�7�F��@�����$\ۈl'+�Џ�׫�Œ��b1O$��HY|�5�KU��mX�lX��6���D"F�33��S�:>1E�{�st�m��/�����(�q�;��|-'N����lۡf�8+�]�WYPZa�a��f�����<p۶l�JWo�N]==:��>2(M6,J�P��Ё��e��<��?B�WЍ�n��p?YPˍ�����2���%l�t��CN�����ZιL�F�G�*%�(���(䨫����"#���<65I�kW�m�����k�|5��WJ��,�yXD�T�u��gT��u�k>�*�#o辰C�x5�~c��ӕ�-7юk�K&w�5t��Я^|�N��7��O��|�p�Ǟy��z���.	8
�Y)(`�����i�A�N���Hg�m�nÓM�&�������oP�����9`�I=�^y�u�HJ8��L�炨hS#[���� xx�6l�@7�t��������޽���ߧ|P�&���^����2����yZ�c�=~���g8��®��o�+�q�z��*:�(R�G��s��Q���Ip�ю�o�n���z�IyF�,Y����Ϻ�
�����vY�󼈯l4+��8�����H\�/O�kMCqdl��?00��RvH�,�)�mu7Mb �A1X��;@�*��Je&/��ۯ�F���Eq�/��S��x��q�:v���	��>��p��I�٨p�n(Э
c��/��l�?�'���������j��2q��g����Q��lO�%�!\�9���5�u@b �{I�K�I|}����쌙d���4�;�;��.��x/����n�$�~��4t:�C-A8�-��ٚ�F�L5��ԏ|�Y�@Ws�4��>C,��]�����O���8��������9)��2T/�;Sb��ީ���2�$���a�x�x�ܮ���*C=J ��s�R�d��.�)�e%�杂� E���)�Ж��R$��=35K��M��4�8@�_z����犔�-���ڼc;ٽy��6x17	q�C���(�;TB�Ay��!�E��	�jo��
]����Y��8�2����4zѮ�d�S]I������U�����J�Yw?dT��o�+bbQe�����4{�O��Ł\���<��ֻ4z���b=m��z^��VNO����\oH�ѕʒS�Sy�$�J���(�x���B3��,�A��m[��T�W��E���8���W��ӎ뮡t:#@��̌�P�]lB�#��j��Y����X ��?
ƞ������=;Fw�{�SV� �k*�E���v�t�'�i���f�i��j���mf� ����2�<�t�1�`ɴ ���Y���;���_��9P��O�:�zh7��ERP]�w1k�N�
�{x�WE��Y�g�b7��@E3��&iޙ3���]Lg�˭](���vi�e�{�5SФ�ku���I��_���JqG�B�P[�a2�:��>���U�� �_W�Y  7���n8&h"����M���ɮka�8M7��5NE���w�Ҵ�m��ϊh��'���+��Ā�j0;x��L b��5��@��݋̮�/K�m��(�_���k�҆�WP��'[�&�`[1ʂ�R��K��Eu��2�6�ݫo����,UE<�Auϡ� 78� �q?(\���I���������t�6��diʩRe�J�=�3�9��}=5dh���b���������_��T��8�'�J�W���\�૾���4�$�rt��W�M�\C/��"�����MM�Xq��׮��u�h����w�?� l���{ҩ9uW2J���&�x!�=����P��ZO��7�z�~���$`��?��t���2F@QX1�Jx�rN~�J|�T�V��Yo�ؙ��lPoo7M����K֭��Hv=����o��]Y��{jSt�mx �*-%��w?p��;. c�j�9B{�������&>/B��G�HB�|n������Э��FO�� ���mWh�Ê������KC�AP@�2��t���(�\䄠�s@388$4*��f���,�U���[�����'ߗ��,�]Vm�^b�L���u�\�\�Vf��4o[�·�L-Pj}�dm+�{�u5�)]��.�Q^(�� �{��Q�%n/z���ǢBO �5v����1{��
$X�߃�����*�1`��G������tZ)7�= ������v��L���E�=i� *կڶ����Ɠ�_Y�e�0y�e"):��=:~����#��ܺ�V^������p�� wǀ�������ꔴ���d���Q:�@��g����<�߾�V�P3�b�Fnš(��  RE���U��@�GѦ�䤢�솝eGk_�B&G�'N��#�hz|��ɔ�I�ɸ��=��#���Z��ʝnϾ}d�Ҕ/t���i��4]}�v����5�,ZEݠv�gPD��=�~�=��	=���	��Z�<u��}�Y������_78�-ߝSn�M�XDE�܄��b�Z�(�^���6�^��b@1\��%���o~�����V���҂N�,_�?+���a`]b �۝���|�^��.������;�~��U��WkR�qkfQH���'}�^z�E۳x$���҂�Vϳ�$���M������(|�+�����BDM�ה�6�a��MhJ<��z������K%�UyKVr�-֖J�,�]^m�^BM܅���-����\5�Z02H(�K����lFBHxjZg�ғ��C�[����7y!��⹦�<j�*�*� �v�����,���H�o��l+�z��F69Tp�T�-Y#}8d��a0�m���pdHP��i ���ܪH�h5˥ ����Th�R����aX@:�eG�w)�H�1HU�e�epﬕ���=���0��J���|��P`(q�UW���cҗ1�����2��UԺ� �MqY��w,��Vpy�Y�2�D�`��y���Z�.2T7�p�]� 8|�����QBFw��dU�J��OQ���V^s%Mzܯ���ܦO�t�\��U�Vp�sl�cEI��*Ś�b~rf���NG��M��?"j�vl����g�zi�^4�5 ���p�����)���0"�l���˸��t�l��]_:C9�78����������k�(�9�5�>�h��"�2iџ���b��h况���}e��3�R��m������q�
t:�s���yo�V!�]�9l��qo��1ھ�*Z�~=�=.;=�����Ǿ�n����_���wm�������/	�v���}�f�$+\:Z��ȜkÓi�7���?�'�XE����y�d�T;���+]�l��&fi�7���,=��Ӵ}�U43>%��^}����V���<E@�@!'�Ʃ�c�s�0|�����o�y�f
�v�Z�w�Q\��|�uی%��i�3�
�|y�\Ϭ�v<Rʥ����3�6���^��5��~�Щs�[L���w���̝�0�bT�4a�фӥ��V�c'�1�l6�\<ϔ�u`.��|LHǙ�����>K�B���m-�wk���3���?	�vs�6�J$l����D�N�7�^R�V�p��@e�_n����h�w�k2�ʈA� �|1	��a���>�m�\�ۚL(Kd,¼�0�l��j�������|e�~Ӈk���(��|�y��Y�H�q�����, ��p#�p���d$��t���>����}{���n�Y�V,�1Qc! ���k��/�$��|,�0C�|j�F�+b���������믻Q��P=?� /À��R�?����_��G�;��_w��[)֗��y���q���Ak(��5F����*�8/<�	�IY�"�F����u������Ӂ�{iӵWS��U,P�'O�|����
Gs�
ݾ�)p��Nd�@�HD�d�?��24 ��8m^E�u�tr�!qsK����z�I���x�� 0Gp@��@��b�
#C�%c��L_��UJFSm*'�I�����6�4�����ŝ�&���#����Ѫ�+��o��}�;��K/��4��;n��>����=��?�3:u�4����t�͔���������/�Qя�����F~�����t����$����辝��k��F?��O��n�`�mTB����i�T�{��h�����>L3�@��O�ǿ�_G=�����>� ��"%�6�}�W�dvo��F�v�z��Wt�����W�� T��)
Q�7�TU|�/�(�����G�� �1��� �<��������v	�5F<�+��W��^2f
�z
�:�y�L��)�^�/��ܶx/����
3����D�����haw�p3�[���������~�X ��G{�CNN-޴(>�[St�Ѹ]�f>vT�"�A�M-�n�٘"y������/Ej��/�Pr�I���;�<r=;=.�R��nͷ��X��,3� �5���{W2��Z"�Ȇ�5u>߁�)TKe3��� (e �`��c�]�&��o�C	p��K�ʤhŖM�~�FQQ�a����� ��-��dM�#c���zե���;�֠B"-� �La�*�K��'�ٓ')�b�
kGh���4�v5u���a =S����\2y�68
�0�^�^36|��9��u��g�l��F��T������t����E��o����p����g�N%hd�z^���L�2���>''�fܖk=��偭%��ɮ��9!ЁTݩ'�瞗,7��`_?=������?&Yܧ~�3����K�7n���LM�Iŏ�G�f�6������{y��顇�����o�8GSS�41v�n��fڼe=��3t��~ھ�j~�C�����o�֮���,�qd�*�GJ���ྏ?H���7hU��R5���stl�~*PlU`�,z�|��y�u�]1*ٹs'�~�mQQH����t��n����h��#p��4)��Z��P{`I� �� ������i���O��6�D9}���,P���A/�5���d��N[gA�?�fvB%��u�Y��S��ƃ�b/����x/�f�'���-�.@�;���h���=�����U�۹����6��Cr8�z}��'�! 懩1h[$�{g��M,��f 	��Y�A���5�A�o��]�|���)8�GFbqZ��
u�#,��TZK���� �?A]p����΄��1��M�؞��G#���͛6����аd����֦��J�h��oPc�H}�<�UJKe讝��,@g�Ju^H�Aa:�a�� RJ|Ȗ�\j��DL�uV����	�ON�q��Dd���_����<E�	Z��Z����y�:}��YE�켛���tE�����)�(�N˵"0�(-6��ZU�5Ҍ	=#�?g�(M=A���Mݙ.Jg2t��MB�=A��y���'�WȞy��W
�v����T�u��J^z����n��Њ��W�c��,����K�==`}��*���+WIvt�����b�q��;�p q����wб���o��]]�m��422B7n���G�_�\�<7n�/�Odv��~�mڳg��C���@�9���}�s�"�v��!D�� ԏ��r�J�Kg�Or u�V��)��S�n�mi���*$��o����׾F��J��:�dvI��NR��\Q���J��H3�t��xm-1���3�*�
|�c�+;��}�8'ǭJ��.��Ep�O�3�Cz�#o���33�E\�L��"�����T\�@ ���e�{��e�{	�Z�*�T �щ��D� /Xl�7���Og%�e�8��
+��L�uR"�c�3plq"�%��z�y�~��W��Fv���;ߧtk�ZE�@���0�5'��d+�_RE[ш'2�a�ؙcu�aѬ�+q��q�EF�JQ
��Z�VZ�!�,>gdw|���Z�3��'Ȅ�"�Ы5[r��"?dX]W�L&%�E��pm�����+$�H;B�������7m�亮������g�j�*��N�$@Q$5$%���F2J�Mی��a������6�=#��I����j���4W���B�[֒����s�}�yxDeVea�d!��Y���ϟ�w޽��j������2�M�a@��DL����9*�VpTj0 D�%�	�¸h��ҏ�J��-�򇂣j�I�d��y�Y��s�5��4�?L�S��{`��L���8CWΝ���Eq�d�?�}���x�H�ǦZ�*�[<n+u��E
N;��Y����`��{�.�ߦ���c�:eri��p�q�-�9��4e3�*6h��Psz���*���E���}��Ƚ4<�GY���ţX�����ͣG��;ǩ�M����p,%t�<�����4u�q�B�|��}�g/R��8�Iĳ����K��pںo�կ	�A&I��4�}��R����b��������qi���Р�Ø��nh�<ϖ9G@X[�j�8��,-�SO<F>o�*|�!������R�788L_���D�� ���N'�������>,��_��Dgx�#b��+/�}��G}�~��_�G|�^~�5:���=�}S��ӽw������¼�W��)���d>�_���&���O��g?M_������R,pDi��_���cO���"j 1��fQ� ��y��D���O�������f�E���t�7& ��YC�����<l��f0R��J6T�3�BM���WA<��"�P;�<��56>.� ��*|��]O����K�v-�n���(Q=��bi���$�˕�l ���|��X�E��2�ij����>�H��ŉ5���ƹ���)�l٨��c�K�1s彶p�}2�xѓ�k�1ϙ�s�Z��[�@(gf�n���'^�ᘧ ����oX�K�h�����<����Ƚ�~q����4ٝ�z�w5I!�"_��J��
���Ka�����S�3
'쎿�aDռf3]�Z&HX��9}Z&IY�b�^,;�kd�Ls47���J��)���?���ݾs�,~����&��`���H�V�R�i@��R-S��
�Td�uù	��_w�|=	�	Z�_�_z�!�& ;�ia�PHe���͕]8s��h�d&��|���*�/�|���*���>)�Ă�;8u����30�t�8M�,0��hdl�f._�X��h1�jPw`�7KRñ$Z^�2M�o��X�}��M[��M��ѩc�����t��
�mf�mQ�rev�.,�(��ٮ8�
<_�e�GG4�hqeY���|�rr[�%���R��T�ƹA6��>��d��f��˝�k�E�#n���b�SK�r�ke�.8v*��}�\e�a�9���W�R�u��]{Ŭ�Y��X���(M@=Z�/��"-//���b�����+���ǟ��~���������o҉'�>��'�G?�1]�pA����в��<!����t:+�{�L���8����F���'���O��y#�ך��������P�Y�jQc@4��S�H+�-=��?}F6S��f��]~M�Ak ����S3vۤ������ϾV��yY�
o ���"ld-���A����q��4�¢�Z�]-:������w��u\�}���Й���Y�w77Q�d-��V8�؊�h��[����+�3�Q���غ�)L�',����� )��(����w�\���[L;f��
)D�Am@!�o�L1_ߪ��j����#.~k�	�B���D��λ��~b-�r�R��u=e�ux����뗯� ��VU�5�{�ݔd��/q\U�g��'8l��7�h>3���V>�\2F[��`w��T�-ӥ�eF�(���$��\#I}���� �R��[�π�Zyb�.�jT��%�(�]>z��MO�Nb�� 9�	�������*V%�M�)'�F?.��Ђ�D��"e}"Ѷ�������s�05S65xV�3Ї�X<�nl�?� �"��Z�R�.�:˳π�Zn��w02 ^���V�^7�A»A�~�W�%��!��s���n��9::Jy����{{��~z�9�����Gz���̙�B_ -�?���H��z��'�|R��
o���o0(O��ؖ��<WU�����Md��/��zH�j��$ml����4{���+�ó'ߥ���aG�\�%�܇����>O�Μ��������~���	��*mC�t���Ҳ���݆j��-��h�"/�h5����E6�N�(LՈE#��7S��/<ߠ��exE���wol�V��b�٬`���X��	e�u��������:e���2�RXG�o�u��*��J@���ٮ��*$�7������K��^�h--��=�vO���S�/�~����-�YYY����P�*mT� 6���R�d�ތ�B30��Z̻*��P�����۶���j�L�X�V�J4��S�����;u�A[��$�L��N>���}W� ��CC�Ӻ΂w#�/E��-JHC:���&>r?��]={��._���SbBѿe��<�5kM)"U	1��0���+� ܩ��pv�&�8M�M���R�����p*G[��hx`���q�[o�s����I �U4���ةw�T����Y�6���R���4{�2m�>��:Ie�L�AE�7΀��\�$ ^-K:6���@稩�*�^��$��-����U�#%k�Ywt�l�ppxAuz!)��������Bfn��>���l(�,}�3��c��ҁ����3�A���@�������*���;w�gh�^e�26:F˼A�����1���*\����::�_����3o���VW�Bg�>A�<IY� ��HT�q����lӧ>�����9�%r)�P5�@�`Yn���^�!�Ĝp.ꘛK6>�*w5H��xߺU
�2Nzm�3��`���v"fB�Р0������6���6��90�7����w��M�Lz�N`��5Y[�ꈆ��s�AA��#�I��ӭ��JtOl%��Ϻf uEj��<>#�U�t�)���%}���YТ���u��"
��n�Fwv�f
�"�Ij�Ĩ~��ZXm�����(�R]��gܓO}�St��1^�sJŀ��ȯ�5���g����n��S��c]L�!��>6#��R��4n�W1�B�
�x���� eҼ�-�P�X�J���R�^�a�:�U�=���.��^I�7�����E�+x�����SOɱ ΰ��|���*�1�r�<-\��Q����q�0@M��Ry���2�8�g+�ҕR:RfL!�/�NL��Q�\�Q����J0�ٷ�N�~�&N�c0�0�r�~�D	����������������c��D���r^�"��X�2�K��E)L�3�[Et7P�c�K����Y��W��J;T]��ß��wY���b�H4�Y����w|����������V+P��e0�� Lб��؁,,tQ�.�"on@�p���
�R���@�!?�珱���~�r�Yg`�'���~��R���b,�t�gT,)z@__o�бwNP�_��������"ZD���~�{�m�=0E��<�r�k pl��M�ghui�
�+�Q���G�E�-�����~���3{���q�������ewo�jВ�$��FKm�������_�"���4N;��L*!�1�ҥ�52�1H��򕜘�+��a�s|9o��@͉!�W��*�E�G}�}���u��MM�w��;�tj��j�50����	
e�^��<^��`~�|��~�0�W|ވ���5Q���R����9���\��qn-m�d��ZYRU�V��[�9�Ex���wx�k��R]x����\nՔ��/�^�$�Z����ba
�n���Em#�����o��a��z�!�s��jzvN@�_B%<�6, V0��	�|�h�2�X�j"��:%��ڵ��G@%"�>�s����Z���(<�/��f��^�k/�Bu�1|^��@����yQ ��7�k8>6vS��THe@��Z�7�@g��ip|��ǆi�������ru��MMqn��1�=[�o��@!"��~b�+�r�R�����Zތ403�X)3�㵭�@�� �Cq�Lr�/ol���<�Ǉ�bJ�B�/^s��F�._�NC׮P.�_j>�)����҉S�iveQ�����ߋ���;�k� ���hj
��B5���G􉧞���a���
��jeݱ����D�P����D�ڭFM��b �;j�����b3�������?2���y�/i	>�=�<44��ϥj��Ǖ*�K��c#*�@m�y�(4���-F��۾��ʁ�!�q�.���ir����1��s�)�����!�� �X,,fZ]-�����;���������lF��Dp��582V� ɕz�@�L�y�b٘DY�kܛN���5�2[Zu �
�T��_$��fk�!��3Ʈ���;�� ��TT���5��fif��}ح3�n��5L�?a1??/�?@TH#Z%TMk�י(��T��r���DM���?RDB9XY���vM�&	E^���.���E4�ֱ��~�14����D��1e��	w+Q�jR��t�4s�*�L\��V�I�|?��^��2B��2y	wA�U2u��k�%�x�THp��������oP���>H�7���k�����~�k�~�=�ν��L�1�C��rc��F�������ɫ3�M��|NŕU�p�<U�UQ��[^�U >F��S�?C;����c��f.A�z�,Z��i�V�zi�.\�����4{�,�o�B�=�K@ӓ��������N\����Hd��3��ϞW�-[�i||�������[˗������5��rT�O>�v	1��
l�R���Q�j�����O��v����l�BA�/ރ�?�9���]d�ހq�h3��( S�ʾ�3��;��s��>.�HV[u�}��x�e)�/E�n��E۷��|��"Å�	����{玲[�҉��Z����[@kSL�W��(]o��-�]�1�(����Ł�0�����q��v�+©��c�G3�T�M2?1u�з8�KGi%sc��oJZ2�^k��̠��U�(���;����&l!���5i����6�_���Q���>B��]�cу$@���I�ㅜ��M^+���߉�::�k���/*�6D��H;�pn��=#�AF|�n�ECu=�K��ʑ�:���ߕZC�R���f�)5��k�&$��h&���< j�"�x�o1�mb�@q�OrmR�ޮ�
_�	�i��׎Q��J���+��N�"�T�P*�����i�n�|/��
���3��Zb`a3��	�
a�4k��oei�r��T��=q��:~��e�����-�3خ��|^e�F�o�8U\����V���Q9e���=�f ��܄���W._uX;_�6Aׯ^�/|�K4<2H?�y([���>@6�Ơ|l�o��GG��Ϳ��@�订��TPW<���u�|ݧ~S��᳑j����}�_��1�)J71& �h|�gH�a�,3����ù"ʅ�2��߃� �l���{���̌ �i�~�����6rA�=�̈���KO"�`����a����Q��ؾox�Q�>+��Aq~����Pa��`��)7.Z�l�+�����"ݵ� ޖ�F�{3-q奮(�*����$M�~k��'���/*;�u��&���(�I��E�CI������Ŗ���nC
�:a
�1��ڝ�z�w5��f�!R�h=_R�h�n��f&oD"�r36��5K�����I����8�� �R�f{�ߺ㴇��:D+�ͤ�t_m�:��n�~�$��u��h�Ov��TA

���y���JzH�� �>�9x��d��Ϳ���H�s�:-���/������Uh|����!G�	���:�S�X��B�����2�,���&�gU��Q֧��%�2%��2�*����՚җ�>�X*�l�W�j�N�466.૥��3�/��1�h�^���o�X�_"�� ���C��,%�&�xW�'�@"�1��k�7� ���h���U<�R��*���Ңݠ
�N�R����u*�D��vӞBٙ4]>~�ܚG��)js��P,�{Zix��r�*���b�ƶoa@풟�Q����?�x<V�:Ň��Z�L|jp߭V���߭�������)�]�M���y� ��@fr9*s����|~C�ҷ��6MC��\Z���`��$Nvss�t��ò��8����l6�4�Āt�x��l*M��W&&�Z8rr�$-.�P�?K����/�㺸�$�\?�`]ˀ* �A���O�i���.��2򘚜��n*.ุ�(�m�7x�!U�I��N(�[�:��1�ʀ|bi��y��/���E����J'�x�>���|���ͦ�Wv����|����4�g���}�_.-.��Z˧��ݴ\"�"a�Ws��i�p�ۼOpzA��\q�[\Z��&���-#4=9%׋,�(o�gT��w�a7lno&cku�;:����kD�׳f�� ���g꿙�P�n�0c����զ �Y���M��[�C�磺�:J2|���|��� ��8ʓ��OI*�V�H�w�TKm��D�p�}p��?�����~Wk�� 	�.@Gwuqo��z��;�� �&j����)��rȢ����9���kX�L�H¡j�x,�"�޽��~�i��}�]����B-����\�!"�Z�ޢ�Բ�:R '5,28�۷�M�.d���ࠥ�䗖E�H����[�
�j�]��5�M)�����#�J$9������m��"v�t)Evw��K�-�B�L���5˅Y��Re��N	y��i�_���X�ܠ�G�q���sZ%��E2����y�P�� �huy��|��ô?~�?7��'ΒÀ6�a[�s��@��z�[��}�?B�c�H94�,QP��!ɠ��?� ��=�%\�ؠ�)��}���)�4��=c��4���������.��I��.-.
���QlHP�8� )�l>+ g���B�t�Za�$)��):w����H�l�Ҽ]_��C�O��ݳ�Zqf;r���'���E�׈�C�aϞ=��F��ߢ<���Y�~��!�0@q�sV���91��fp�����m�=4��!'� ބ_;s��v���KSER���\�y�a��+/�F8� ����~J��:��x Z��:`�f�n�C��@E-��-��[!"�pn������iЪ��wo�fic���&8[��W��f2���FѲ����->�3굏�� �&jH5bqp¢&���ֶ:�i1�W�uo��RX�d�N#�Q����!��k�N����-z��Oҋ/�H�._�%x�H�b�D���5ŧ��Xz�_+����0��h���J�Z�� ���T-_�["�p�󔲃�\,�έ��/�?�UJe��$�&��y��N���Ha�Ƶ��0�2T���ޥV�P|�n�QZA��ЪW������^~���g���"�L�9�_�+~g:��(a�Y�ё~ڵo7M��H�����X6����	�T�����Ya���)Jf�w=M�BuUxé��d��[GQpK�Uz���}���=��#`���S��Hd�p����x�=�e#299#& �w�}7�{�,��B.3�:y�^|�eѰ�[\�8ŝ;v����ك����; ���wD�Μ=�?�t:�2��p��}��ַ�%�
�ߓ'O��x s8���G?~��y������޵[�e�&c��3@�Z=�㕿�~ N�|_�����-�0R��
�N�s�>}h����
�۲~N2����<��C�
?��6 ���|��iB��r��A�8�i.�	P :��~l|�Lx���k<C�ލ4� �Wx�BC8�A�׫ƨ�o�A�Z�]��7W�3��khѵTv�*��Ū�>��{6Q�B$���YHա�(�?�D�T��M��-�f�X(\hk�X�� �#tB����c�=Fo{�^{�5hH�8Ԫ�P��y�,z>�S��\<���VP�h��Յ�a&`�C���]\�	��V�#�gl>Â�5�t��ݶm[%�W.הL[���dp�7��IZ�������� u@����q*���r��
إN��L���z�Ҥ�JE��0
8��闷��T�6=rR�l��~��X���|Th�b�F���L��5Z%� 
�X� �y�n�z����4<y��y>~�ټ���B	  �q��,I�'S	�l��] �ne ��#j< >poy�t��}�[�e``X&~��ࠄ��r���>ǀ3#잻��k�r �uߘ�����}�1�8q�8=��ct��Ò�G����gX��={�._�J=� }�_0�����/���6x���'�?ӕ�+���}O�؆�DX]1I gd?���O�틈62��K�k�?�3�� �[�l�����$�J�.�-���oz�<v�����/�
#͆ҏޱs'MO^�@U�\t�[����Y@��Ձ���*hb��/Q��@����O���3/��u ���X�`٧�*\�*�3o��ϽӛDxu���Y8R�9B��ׁwP��MԔdU'_��K���]E��ꯛ�3:�\��g��_E[�o��M��Zʛ]�웃V#���������н5V�������ط<�y���q���y*�L/<�[����L侼� 7�&�\��
��d�5 1X�/^�(�w3[	��Ɉ/�Tp�=�v�Itj�y(�
bU��j�*rG8?%�K�	娤�p(��B��|�H��P�3��U"/Q���Ⱦ��~磟|��ryjԚb!�bP�t��@,Ѱ���P>��t���Ǡ��&����-NT8�1���L��T������6` ��$X,A�b���8O����-��*���Y�9��W?3�����Z���%��+�2w���,���b�~��1!�5Šhp���A��%)����sg������m���2F+�p/dL�q�'����9�v�����%�k8�e2y*�����m�,���d��;��c�"�U�{��_)7�1����_���[����A��7������k�.aP���Eش��BK����������L�.��D���^�oݺ�q8���o�ֿ��0��: �i���ǀx~a����/ϔI���-�kGs�����@�V��rO�Ж�;h��Um�ƀb�So�O=�Y*M��s���k����N��#�=439%׀��s��u��.�R�6�<�����%nq�ë����R�H5D̹����������Ґ~����n�걸I}�d����;�s̛ݔ��@�1�	�_����H���:���.~��-�"/��o��]�૵xW�:+��b�V��4�ڝ�z�w��6�wꚤ��I0ٲP�"�n�~���fk�m�?m �������� �mR7�}����*��*�4 cH�a����� ��6ł����J"��č	N]���_�x�&�����O�dO�XRx���Ⱦ1���i���9� ����x���t�i"Y����4�0�a�2R{r{Ł-�k �����bY���ϿB~2A��E�L$�HE�m'A.���e��4qy��d�m����>����}��$(�)��
4��f)w��p�S�9���N�.���N�M%P��W*��ٹOx�?��?�B	�
~���"��Y�� l���[Z^���u�x3��,�,ʘ��0��*���(��K���r||ƭ~�w����#G������|�M��=���O+mQ6�e�56h�N�^1�c *�db�֭���$�}������&�~���཯��ȭ=�������}6��o�ǋ�F6v�����I8ܟ�ܯ+W��CZ�K�3��q��j×���k`�S�g~��m�T�(�(:���7��������j�����G�w���� ��|ؑUR��?�#��U��{�5�z�Ѹ��h�}���$�"�wT��MԪ���������
�MK��ڇ�  L��<R�"�/Z�J��ʕ+��|�$
��TD� 
�\S7�R�4�t�q�k�����R�m�:Nc,MO�a��%�� ��hȆ� ��Cj���Ӑ�T���fu�00@���l:#@�qE��DOWf��-��>���3�I���&F/>_��&��������@sݫ@�$i�t2K�sK��K�Qaj�F���-�����I�����<{�jM��Hy�3B�ܶS��?&��f��9�.�z���t��EZmUi�R���`&��������(%��K�A�������u�r��g���ӧ�Y��N�C�bjvF6Mؠ��~K
a�066F�kW�KY ��������*_O�u�_�@Q�7��M�E�����K/� \\ �O>���_Lk�n�sx��[��O���/-/���yx;�ޱS�O�{��}K������b��=q�$����b���瞣��!-w�T
$�uK�*6�#�'pA�q���+o�FK�Qd���:-�����>J k�(�G���C�s=p`�D�%�$Cy��i�7�rL�6~:^+�d�Lf��P���W�E�#�<Z�M�Ԡ��l+>�榓}TͲU6DͯJ[9,�#KQ�x����J�~f��������aA3��h&eoROEk�/V��fmݾ� "�@2h e!��
�ر��OD�<"Z ���k�D�ָ��@����}��mg�v���B ��jY�[V�
�*�+z�p�*�讦�8�F:���\|dl����dUR_c��Ү�h��$���7Zu���n�2��)���b�t���]�������P#� ���;�OM;N��KG��&��Eڹ�:�����ݔI��]->�?�GϿ�s�D�o"%���⃇� �������k��Ջ����,�ѿs���*���h+�=�hh�V�Jq7-�n�>�}����~�����j�Je���1M|���x C��G�ہ�6_#6O ��v���" _D�� �7�Q]^^����g>�?/3��1��?f���v�ܭ�(n;r���7�|S
�u�yx�w���}��������GyX�5ę<k�&�R���?��@�%�V<���[��V-TG�MT�r�%>�B[��<�[G���.�ϐ�@s��B��-M�Ҷ��y���wMBQAQb
�� ����LuZ )�%D�{���L_��զ h �92~��"�Z��hFJ,j$c�!z����u�����䷩������aa��	057�V����DzLA�oR�F���*�;4%Pgm�n3Ś[���7���P����hެ�<�b�R�~�}�f"�������V`c:��R*0z���>��(��� �b�D_غEx�}y���HA�>u����r;]��3�Y��R\F͎�1�� ���Tb���
}��gDr�lƕb 4 /��R�h��W�F�BH����8v<�4�Y*� }>_�����/��_�e��-L�P��U=QL�c�W����ܒDR�Z1z��G��$��ZԌ+�n������v!&�U�0�&__\»�_���q�5�xT��4��P�6$���lz��g�45{��=9I..�.j0�@���,�e���U�*���ӡ����]�*�aGFi�Gi���"�뫫��ϵ�������h�����Q�>&4�Z��Ϟ��֦*_;�������D�����h�3742�3f�404�7��bkb��gٵ�#u~�?E�Öl���Z4f%�i��=�������>��S2� }��l�GF[\\9>�)��[�*����k�JM��o}���p������� 6��e,Kq�� �Z)���KZ�r�\U�Y'���l5�O?I���eJ�_���{t�7~�}@����h95�q���_��O�:���I�x  ��^��΁s�fQ�L�y���њ|���rzь�/^����)sP
|��H�6�m�Y����_���	�?�>8�ˋ���X�	D�C;,ӌ������B�ל���-���V�P�u0݆B��u����j-�8�޵��5H
x#�F�%H�u��w��&l�x�7?�O�GAi��9�x7Q����rX�uAi���Ex���l?�f v��.�؈��e��e��	O�	��%�Վ�}��D�/8�BT��\���488 7F2��h"( 9���@��f�%��.;�g��� ��;"�+˴s�^I�	W��'�^�����V��ϻuo F���T���u}�Fꂉ�jfQl]��� �_P�leHȎg��c?mg Z�똙�a+A�
o �M�<*/��J�"��� �#7�'�q�;<]��M��	H���1���p�4q�<y����݄M��,�"���7�'�/%�~H�"x]��
�Uɻ)αz����Z�$އ̪c��$,K�r�@$딲���k�Ia�.Ds�8������Y���;��c��R�v�}�Ӟ�;(Ě�,�a包@�	`Zh2-l�24=7K���:���1٨<x��z�P��6v�] /��:g~�'�LQP�V<ݱ���l
(�_�PB����ϢH�+�G�� l��������	pjy�MA�<'k<ʈ��kϿ��Qå��g�n������=�����ǳ��;�������K�u,�{��� �&j�cc@tw=��gv���a%E�;���BY��� �"3�TB�X��Z��?SS��{X�"jd �e��N$`�V�b�Ek�t��/Q�V��?�F� l?��KV�M�j94��r>�ظ�A��ozz\��fD��<`Zp>�F13='`ګ��tS�|�UZ���HR�ϯ� uρ}�[a���5v�7���\~7���|�y�������]w����fc41;G�+||�FN���&�+%j���e��V�|���^�~���L�rQ-?9IÃ�+P�/:�e��zC���~.e�.Q� �b��g �R�U�:ol��*%SqU\�e��� U�V3	��l~V�����ހ�vgm��ZΑ���y�}4��ω;��K/�?}��t��z쑇h��"��= ��t*?�b����Z����[G�|��Yڹ{/}�W>/�cc�JZ�&�iT �}^�\�jR� rg�϶�[4�@<�ϒ[m��̂O�阼~�������M	 qL����ݻw� ���y�<�, �#!vCv�n�lO鳆Q���`	4����y|�-`��o\�ڎj��aC�_���A=����~���*��uO��]n���Ni=���Rn0�𴬕=W�6_�wQ �Q �;-�kZԽ.��ϐ�
u���I��T)��D��
>o�������sn]w�פŮ�Z�	"��)^X\��#
��'�Z*�Q��鴣��(2�4,�N;[ �������6 R4?4�*���� ��VM��-!(0�L�F�ԎGZ�:��K��?�59&Dr���ߕ����j��St��r"IU<鄘cT�uJ1���� Y�sY�x��ʵ�;��k�L�J�j�]�}�%�䀹J�Zy��������������0l��Ì�7#��KT0��V�X����(4��D�[��y��ܛn ca���'����W��_�
�ر���yђ����g,��>�(�q6W9�Y0Nx����(�Μ�c��ۇ?�9rX8�����9,C����pxA��d�8�7�,�z��һ��^�&�NO����s���u�VJ�2r�P����TD�n�����Q����
�i���i�V�fN�߽�"��otW5<���8�����θ[�n��N�[��q��+"�H���tB�ӂ te[䟦x�m`5�N�����h�^,dH��z�ݶ���im���o������DZ�9I[��Rnk�g����"��h�����2	�u��� �Ե�R��8�`�3~v")0���XDn�C���,&��0x���r?L ؉�������SSSR�F�����Zr8g�&XZ��T�ǵ����4�8GO�S
`sf�W[��W�S����2-�.P!�a��8�y����"y��+@�M_��ZO���k�p�Md��/'D�}��OOLҥ+��\o��J�(�`�M1rU����=��`���ߦV�Ǽ��G)ȵ��d%��{+MT�[°�N��Sb.1;q������h��	�Z�a 6�ڔ�AIG@%�Ye��6�k]���
9����K�2KZK���G��t!���η��'Z�1����4�e�z�7i�7 G�z�~���4<4,J����	
�j՚p��1`>� ������+�
Gd�����i��p�q.�� �5��͕�\����*��8�%��>G��݇����'����ܞ�Z�%'=��դϓ���*j>%S9�l\�~M����&ys�g\�%T7�T��bXT�5d3�_+�B��<�J;���"h[Z<��+d�Z�ϙ
\t�O��r�r���J[o��)�3-�P�*�ȥ!��P�	��茖?�:�����ӟ�,�z�(��u���zH��oܲ)��pM���YW<�f�碥�5i�I���X���u׾Xjo��Q�%�L'����)�x7Q��n����"�"$�M >����!��0p� ��z�t$5j+�PImv#l�Zw�� GҺ��HU�09��`�00�0�6Ⱦ��GDN�����\���k>�N�G|"Ȑ�2Z����k���������2Ē���>���K�h�j�Z�p���&8͸6^;���M�Os�2�"�� ��P�I2pŗ�e׈�W���@�e�3�ڷ����Ύ'��2�@�Rn�4( ��;�O�� 	� e5�2��̛	7Ƌfҡ���*�w0���@?��� K�P�� �O���I��z�lk4��l�h[K�6�D�����?������勗�ҥK411!���j�*�&�����F��]�v��� 
�1�MS�֚��u H��p�[���&���8PJ5~ʫ%r9B}���5���w��Eo0�oika�Uks��5�VB޵�m�ݸ���)%�my�3�m�~����^��� �T2u&���ѝ�zwt5�&
�Q�bKEW%�����@[w���j�6E��ݘ�V�0@�/9!@@1�dLd�8���'���D�Pl�`���2"�yf��E�Ekp�k���ij���Yg4�G���]| ���emL�4{�1��܌��}}m�#ÔH%��#�*�b���J�V�a���0����p}=�J�"��-�L�g��l���}T�����L�GE�:,7t�C4YYu��T~��]F��O����Q�Y��U�(^�9�T"Ii��l�=�0��%)���e�C ��h�A};f���z��ղo�tݿЋ�5;힥��ĬCG��������������k׮w�
�Y%c��{y.����S�#��['��Lƞ�J#��D9$N*�$�Z�w[�O�V���%ʌ��M꬘2� ��� ~^�?��?H���)��j���z �H�����dã��G˾��b[�,n?�a�n8~Hg��돳|��u`�P�L[������Ud�z:�wV��M��l�n,�c!A���:�^�U��nX[��$i�$|�E�^c߉��P�m���T,��c��~&B�j�6L�[�l&���*�:����p��R�Q5`�hn�z:��Z��� -.�
�=��'�Ts��BV����� ���7��Gv2���V;7{�f4�-l <D6�=����$�Tk�ܧy�}� �x.M�-Qs���2��h�ZP�1��zSQ1s�Z��M(jI�sAK@:l_|(�D
�._�&J���A�Z!�8�<��Y��R�� 9�<�	n=�f[Ү���?�L���(� V=����BQR��x߁��:��{	0D�b"�Σ��f�*�Jw����x�)���d,b�TʫTa0�d�멅9��Skn��K�2���Z�lK���l:���F�vlWT
O���G�����&���f�$&���Aq��Co*��Ԡ^�l�����F�6��lMe��������9�X�j5�<�� ���n�D:͓{#T�d�toU?;N�Cm��R�+�ʛ�~�	CTѤ�ZZ��fME�� �V����_e>_��v[w״P��Ɖ��.;,�g���lx|�u�1Sɔ���wp�{gк�a;&Z�0 7��\FI�����J�e�8ra��C�YS�:^ ��0��~��^�b	z�'E������_�z��Y���+il6�Ԁ6�_(�A��^�)�u2�
YR�mY��o߶�-�sY��z���)J���v��D�Q(��t�O� ��lŭ� �"�����,^��Z�^&��8u8�����"����E��@��"e�����6@v���kr��u#ōH�j���Y��R	�2�����t")�㎫o�O���\FG��N��KK�OK!c���{�+��ζ�#Sios������Z�z�[7+��&�5�K���������vGqX=�������������y�}U�.�cA[Y��>wC\���[d�+ �\�7'-��B	�_C6	z^ �3�()������yiV[���(��}����<%mUH	�k�\��^�`���I��%p���T�jPUiԪ2��\�����Z?CaPu؀�94k��v,W ����׊p4��,U��M4��i���W�Ǧ��k�|Z��#��6L�bԂ�ژ
����Rh�|��W�z��TY�s�Q�Us<�P�������&��}�Nh����&w�ߜ��|�Y��g$����Q�?}���\���mG2S2'�"���vw`������N6[��Ҥ����D8���/���7��Cp a]k�z�#Y�o���#A�C���u ������V��R�k݁�M^OJ�|���}�vI#��	z�0@���d�;�WK[T�("�J���#`*��I����<T���i0��`�5����jvt�0˒��Al]Eo�,]X���R���RS�+λ��p;�S&%8�eC�~3�	�aX�;��	?GR�Bٵ��Qe�}��h�oI1(�y@�M)��Z���[�AU�����5i~و�^ksu���G��Q?[
�n��h$Sm�� F`ߔ�Z6}����e���8���f� �����ܤ��s�1 m���}9���b�|������JV������ukfa�|��Y~�y��9� Ƶ�!��k�OѴf��u��
�?��C	���3�ЮW�
��q�,�����}�m�����nG�{�h�F��@_l��x�d�l=���/�?sc�_*ʄ�.��/�}J�IwYdm�����n��`����.f�n����f�e�H`�3��Xh�[��$r��DQl�������91G��e3y�������{��ywˠa��)E,��elX�ng��!_��E.I"XɄv�j*U�u�V�l���2g���}>����>��Y�sD�k|V�}�0�-��N��u��"E*��&��R����m����!-a���L��D�`�N[���O�wD�m]�����W͍|��Im�cVoκ��n�t�2P�������&SI)�����B��C�Ռ���9��BAd�@M	x<�-���UJe�a����z֚��XF�����ٳ�N�:AY����d�AU�`@F� ���O�y<�XI� � Wъ�/,𵺊��[�5��8G�!�3f�O����F�����7����;��*"��Z�v/HtG���dm��-�Ng2���²��ו����=���7�ھ�`e�ͨ < a@�|N @�F�>80���,z5�fA����D��8./�W����j��&i�/�]Q�V����K�#ǰT���C�wwDO�v�e;�,i�d��д"�>KQ>����b���� I3���mk�v��v�ݝm7.� 3���puE���<JQH]	�XT+�J4[E�aG���d�T��L[Ʃ\.����U�J��ۈ�Bk��x�"W�����P���RP����$����ݦ������� 	����P��;!�E7���� ��47��������䩓�)3�k���U 0Д�݊S�B��1��I9	�d�R	*a�5�t�lY�d(�FZ�4���1����"��s��yv7ӷb:�)T����5Ĩ�Ĵb�M�����_�GQԚ�����=�:7�� (p�m�5�Nl�s�m7����+��kS/J~'���L����w��9N3wP�UJV,oSi�TUR� �C.~k�FM1���ȵ8�7=�[�x?�<�pv5�&ެ�|m-�%�jM�L��.�k��`r��t���Ēz�2E&"$@�兯�T2L6���v�DP��_��� ���Ǐ�&$xð��]��+W���u��]�tI �r��x�3H�5A�V,r��EAd\?�<�
�q��W�t��h���!ƀp`x�⩤p�G������`�4��t�>�NR;�ؾe��[D�:�q|e��M�SF�դ�i�__��2�t6�/��v�0Phi,xp�G����e�� ~	4�@q���4n-I��QD�4��F\�.�똋n�1��-�D��_��^�M �'�vd��k+�ƿӦ	��m7�!%&�yZ_���'&�ҥ��,�����1h��9�n]4��r$� �~I!����Ҫ���kuJ��o����'jؐ)�����(	��(0������O6�Q����Yb�a+�v�֔�f�aC�b���Ѫ<�`���Z䚢W��ڨ�8���P�^��q����"��j�5�+��~�"�z��ѳ�a�o�/�}�5-��f2hvW�iBK�Y��=�j?,�5|��̉	��2]�헹�W
0���8�ɭx7Y��ē���E���H;@ �iA��{_-�;7�'*�3Z$f��B�.�[u<[HDЍ��m,��.^�K�ظ���������VVhnvF�Z^S>�PX��XAC����Q��u%����4wo~�@֪
KA ��)�@�h�g7��P�\�}���jŹtZ��������#����I3'�k	`�����jl'��$������(b cf�o
���&1)�r"+qC嶊됸�\/U~����k�<���rFߺ-��
>��H[��z-��m���Դ�D��3����a �lea+���۔±����H�WViqv�|�BM��@QA(��F+�d2-����>#C愊��ϯiOc��*4_xN�4�z��RL��Q��mH')t,u�D���<���.@��{ڱ����� ���ɨ�t��z��� �&k��c��N���<EZ�@�_��6_k;�x��H�K�.o��fY���'�퉔D.Ҽ8"��h."����2qET^|�%�Z���)���p	��jQ*�������܂\��/�-����j
�e7��/<L)���,"�MQ
2l$��),
  ��[�2��)頦Q��t�P�r4� h�� ��*5[�P�$&�#���~�h�2����؏Q�?����5�]N�W�h"�81Kthu�����a������&P������@�/��Q��6p��<K%����v�+-rdA��p/k���EA\��wui���RM���X&C� �B�es�̙g�q=�5�f��<��:]Ű�Fx�<��*6 }�}*k��6��պ��j=�84�`i��v��A����
�4��@�X̙H�Ԕk���{�������X����J�j��k=���Z___��w����G?�����LTOh:��HY*����#��LZ�8�4/�p��X�y��%�"��u�p�B��  |�|Eh��i����y
�Gyqs�4ZX���1P)w4S���di1���u��|��@$PZ��3�p��UKE�`� p�]X)�!�C�:���� ����D,!������������@�
.pv�P̨/��_~�k��y��������|�W�h�v�3�VC]�^X�3�n��`���YCF!����wo�o�snw�S^�uC^iI��SBu��u��M�/��~�g�4�'��7����@��c�?�c��[� �DJ�zP��o��ۛ@s�j���F��G�g�n���%��� }h M��tZ����Bt��56���Qqe�At�C��4��������/h����M����_�����>L��h�����y�x7Ys�8���GM�>��I����Xx6%]�7��7��Rſ�ڎD�p���qn� ����� �ۢ^��)���H9z���0��a_0^�-�*��3ܝ��Ha
U��ƛI��Uu�g��?0(ڤ�v좯}�kᙜ�T:�:<6:J�BA���3St�(��ͫ:�Z�}��.3SD��e�?[daE�6z�)ЖYNؘ�J%2�'��G�X�Eu�3�!^Ρ��NE����Ȧ�	�Z�P/��S�8��".�
J�BCD��K��[YZ��uB����u���T,k���K��}f�U*5y]�_�{0F�u���2�p�k>fFR���.�Þ���Hq&��s��;d�L�6� ��D777/�g�;"���b�\,6$����$<�z�J)Yu~��8(��s���"�R<n�	�!�8��+劌�����I ���R�0�&�D���s�J����;yodh�%�y7r�[��l��ߥh�ͫ�0E�-4,����U@+�㦛R�D6=J�#�1�����.!<qQ�Ӻ��t�v��N�����h~~��.���ME�#�%=��]��RF�!
�#ײY�:����:��[
�e���u�M�;[G����cW���dSie���y�;y *�`������������e5~��̗x�A�pu��!\3�q_���� �^ʜ�wnd�S+:�7���2j��s�sCP�f���Fv
R�F3�{��9�g�j�_�F;�D�Yk.�D�`�6�	Ԛ��F*�vD�q.��SUm�M �P�А�{��Z���wV��M� 7�����:����u��}�<�(�j��lO˒5o]em&J TL�X��������/���.���┘��Q����[��C^����9��nzMO;��h3b �/����JC��/�Q/�X�NFT+�r�s1�@�u�n�:�"\����`-�Lƥ�	���fE�?�W�7�^(䕰>��6+pD3������9�";w��-t��%��B� ��rX��OX_���ò}�0,E��QxFj�R��S�G��	�~L�HY�� �������ih�a�������_������@�C����2�w��-c�r�x�oFp��p�Kp�K�&,+ �^���P�n,�����e�ys�Υ�l~����{���S$d�ߋ!,�UІ�bN��� �lblzM�����/�c �U�����Ժ�Bs�M��MԾ{���V}��13�:�t����aos����� 4*�&������mɶq?+����L&S��9v�BÝ�z�w����6���Zv��\o-�R���qV�Y��v�(�w�4���ldǯ�jUE��j��ٟ�S�-"���(> ���¼DL*��
`�?8�EU�����y��V��'˼�fe���(��ݱآr^��ͅ�5�����Ê~A�6h��I)+p�s�_G�R��,���u��r�C��M �4DĚ5 �$�����O��ھ��JEq�����1�]ՆD"I�sK�����h��JY)�+S�7��ʦr45u��5@F�tqn^��._</�O��P��eT"��"Z�� �N��$ ���U�����l�_��cj�-���������;v�҃�=pG��N���(�5^/�p��2�|�����,@x.S���8(1(��PX�l&T���F^S��7���������S��l+T��x=�fKU�H� _m$ ��4eG����l��Zۡ������Kq#�k�!3���uc
�a'��؅��h�{�q36��j��F�=?ٍ�EÊ���f���H.�D�h����^�sZ�n����?Wc0�lI����!Փ��5���Np5���H����[Ey��(�}H�MS���;NK�+�sc	��@Wo��eUtz[�l���w <(�{ߓ��BpH=7�� #t]�^m�(j���N��s �U"�q^Dx}�9U�:"^��"�-� �b^)��R)J�� �U驧����]�>E�rY� (9��G�GD�^Q_D㧦'��Y覧�S2�����EZ\Z��G�l(���7^��^zA>ׄH�<@�<�Yz��[��s��g��󵯖�$
]b�� �b���?��d��=��)�)����"���%9/D������"G�O�45i��@�U�B"� u�c��Y���1PrY�8�!�;�����h8��bQ�[�a��� ���pP,ʣ%��*�]</�Vk�i�^[���xTi�@�������Ȧ��p�4[O�yc��`5���r�ղq��Sy+��/r�΋���HZkkw�0�Ril�B�pgv�Ǽ� �&kHqoݲ�%�%'%v�1ő��j�Ԍ�߼*����t�dM$�[���Uؠ���01��h����#6��Ht�\�Y$6�m�5�ʑu���Z��:��L:��������Z�_�]K�A�`�b�pn��ooX�V-Q�ZՑ'[�r� ��iM)~��ʒJ�7/R\���&U��d��V[��)��D��k���������Lb��س����lfS6������r���Q�4[��'b�*i_ ��g\_X����������������{�.mi�������կ~��|s�$W+r� �'�=A���5�P�H�y�P.Ri�ST~)�J$�)�r,�W�t��9������:�ܹS�=x���'O��_~����E�>Lː�[^f�9�?�@��<!�Ʉ+׀{x�]w�u"��>D�Z.љS�҃>H���!{���7�A=���s�7/����>�,-p��\d��y��Z��&�Rw���k��&����qq������3�A޻w�����?��%�{ߑ#ܧôR�ԑ�n��hT6� ���VU�~DL1��&�UvĒ=�<����Y��ˊ�s��_� AW��*�}(H�����M[�~�t�pk�A���y<c���T }��޴��k�@�"�=G��
#�.߻ h�e*�X��a�s 1�/�߉����Y�	=�pf���P<����kU��@��58�xV�)RLe"6�ź����Zri%K�x�uOI��P�i;a]��e1'�Obn ��h$�zEM�H�(��=��E�Aq�����J�s���G���l��A�(���%a<�`ҝ�zwr�5<��@&FE(� qmϣ^�p�h���.~F�Z�H�c3�	�V�`nS lC�)���"3�k�!e�,����t=x�p�ӛ�4���h��f䘂@�pnbq���כb8��U����Om#ȩ�P&ᐨ�ZJ��H�J�������}�M�2 �G*,,�$NM"e�e����m7]�v����o�k�������+_�
����ϟ��G�k3t�����o��޽[�$���_��[�қo�I���w������0�g	��H-�3�8��tB4�㉘�G�����R�
oP������~���>)P{�嗥O�������{�[>��/��F�Jr�����|�À�<=��c�����I��o�kJ������x:�	���/����ٿWV�|��X�~��&&&�?��\��r�^������"��ߤ'�ܧ�����fK���.�����9
�Z����v��Q:R�+����#�����n��	Eϙ�Ȫ4�.�(����z��m�iU�.B`��:Տe��k����00q��x���VEmxma�����z�;�� �&k�Y�o٢�b!�5֖���6�Q���%#H�Ac	�P[���#@�
��Z]R��:4�	�D�~2!�t�7B!��*��m���*����Y�l����0�ͥ�H) @��Q_-���>����ؔ���1٠v$�Hm�2���F���lc}ȌY�Zv �e~�ĥ�����{�҅sq�HG��L�����K�/ѫ��@���_3O�F��)Q��H?}�{t��i}�W��_�Wt��y�e����OJD�c�T.zBIx���infZ6 � ]@����+����,��������p��7��u�خ,-���w\��b����!���۷ї��E�?�7_M������ߧ����[G� `5��|���7��k��0G�y������~�ZY��Hs�U��<(c��.J����E����W�Aub�����20�q?�Q��p�1���!N�ߦ��ψ���<k���t=�G�<�m�ʗﱔ9a� yzS�E���^C����,c2�Żng0��V�5�@P�k^�Z��9Ft�%C�ȯ6�����z�w���@`
���up�x��o&�h�m�D��n#�;H�#m�H1"�**�"5���ҟ��������D���,�C�����m�i8�J�H�����C��s"3�2ر6�J�������ʴ����<��k���y��3ٴDS�?΋���_:K�+�!Gz~~VT.]�(���ߖ����0�)ߗ�'R�R��G!"��&.��2---H�����򙈆��w��M�0�I�T��t�={���F�T�������a9�#G�o��t��i����_�uH)�\�[o�%�E�P0r9������"=��/��?�Ez��W�����B�%B<=5+�T��>Ϋ��G���$��(%�����!z�W��W_�c?��S�I��yo��}�U�=���/����[�T�������]��h?7��n5���s�ߡ:�c3iٮX��)��>�V�A3*7Q=s*�CںRΤ�q~�%�N�%~�M(���\8�JO�cc��Q��^����Q�0*�ug2�r���(�O��#����Z�n���W�F���/��Ņ%^��P�@�u��g�=���+�s��U�r�Br"2H� �� ��%YV�l�Z�0�-Y=�eO{~�g-��L{�c�m+��-��$�
��"	"�ȩ��U��^�����9�[�Q��:X�
��瞰�>�۟1�/�4�Q{�	m�%.<�Ҷ<��9�o�0YAD��1h�uTJM���VSf<�=�#76�T���˫o�)VXo�݉Mv��\��?~=�fg����BT|Q P2a�vydV1��f����>.�&�����3�R0�c�	NlF�F�-�ǌ��������|��[�����[�%:	1�[���p��e�Rx>ӎ�^`�9��8���N]L��x4�"�y�?2*�^�x�J|�%ú��в Għ��`t6��J�p�����D�(�j�U�KW��j׎��ꫯf�؋۞W���Z�hm�\�e;Z�����h�UT����Ԧ���X�T�Z���|��������� e �V��J���������Ƴ���`����N�m��� ��� ��r���~�z���{٬�-[�6m�Z=��6Y��nR#�#j����b��>�����i!m�Sյ5����$�"�n��&������Cr����)O�߷��M�N�8��X��r��}^���ׁ�҆��Du��$
쟕��+ 0�o��`%\���&�x�ԼF�h�"��1-�q���T�������X�q `�k��=�=y�	�|(�k�;�U9y~px��6e5�aV>�3��;{G&��Nh�b0��eү��k��׌$/�#9Z���5��-��HAc-��^� PT��,�;��A���lkؒ���Z��Lp�8�bތ���"��y��q���=q�ʸ؂��9�= D��:�_�b�f�,�����1s>{,��ģ����Y��}׎o8��_&�A]D�J����㜉1̐����./M2��---��ղ����)S��+���	S��2��"r��LZ\@X[��c��7[0Ir�5�C�*��|Bah���j���:1�ɠ��,����5S�U���g����n��sv��y:6�Q��dI\�������"�c�dDY9:E���p8Y(brk�h��&7�lM��766�D�g{�-��5G���K2A�e1D0+��	���6l�R����J���]�|9�N	v�5<2��eb` �����(��\�ջX����;��������jhhd}-_��׆�O�>���r#� �Ŭ�Y�c1sf'3�e2��'�V�x�I>���j�5�rr��13ԇ#i�u[�U����s;,�e��Ԁ�Cǃ<�-dh{!]X�t�z������ ۋt�3fLg]Ⳏ���|�����u���]�J��������x�!&yvu:i�;!���^�cA_�Д넻I��s�ң7bwm���Y���٠�2�`A!�Ƹ� W�0�$�V�?�M ���x���,�W���aLt	%lЀVk�mr��9,҆���LՏ�x�*�ye�^bE[�$X1?vR�D o\4�qq���r��zŮ���E	�_���y|2�v{4PȦ��~ �l"��#R��5������	�G4@���߃5��K&��1lVe� ݮ͖����2n�a�����;��8� t�c��H�(g��Y��!���#�hӫ,� �yU���4�LS��p�jl��C����������|�r��~��T���C:tH-Y�������{�ڵ&
?��� � v.\��VWo����&�X��Ɨ��+ � ��Y�Nuu�U^��5� �v��E�4�Ψ;�[͙3O-X����c����5!��F�U߀����}�ǅ-����t��5��P��}d���^���o��V���.�^��u�i�
u� 5���r�`�p��7��fur����{���S�t�l��z��D�����\�gD�n,I��f\L�=��U~v-kwm&��U���������	3�٭r�n���)�	p60�}%㵋�r�&&��[1���^ֵ���X��w�\���E�-q�q�g��v���h�p<u5#��(}*/��v�bw�oe
�^j�a�XP_WH�,��O�/V*uT��8F�fD���V؂�*�!�[i�ł-b�Sì"ȋ:�$2@gȂ39@����֙Ŵ�$��|�������S����
�o����*�4��a'�C�' y����TѬ�v����jȄU�^��_�Vdu�Z�[�N��!�[	��+&���n��Ѯ����l�Eo��?d�����9�"XRX��#@,������������pLX�t�M�9F����2` �)�`�4�|.8,y��`�~��h�|�J ��Y3Y_����&�#,�jjjQ�5�B�m-�8�:����&�:R:���:_�x	��64&�f���lr���E��h��=���, y@���[�5,0��_���Ԧ�&s	� ��\S��`W�� ���`S*�͝���F�ۤ)����QʒIjyW<�++q���v�u�7�g��Ar,1�I<��p+�~�d���w5��[�&��.v��c4�p\��������d��b8�A�����*��e
�^b�:�:iM���V��F��uD)'t���+�2�:'����-�+e�8ǵ,�Y�W>�·��~�n��#�}<B6�q�2ZM
�e�+�Wy����Z����W�9^e���.��O�=�=���u&̘z0M��>��_꩔�i|��@0<ad�J%8`�!b]��Ⱦ�!�/oI��u�r6@�o��	�wmZb��xze��}���������V�F
�<���k�x�~`�0{�g|Eu{"�F�Ԁ @���^0�q�ܿ��1�FGGҠ�s�`fZ���r&@��\?@-�~�Q�+��X��N����Np�H Z�d ���u|`�h�`V@0 �9���#!!?s���u��E��ǂ��V(h�0���:���#���Ҧ�h�7�\H0��5�Ӭu���1�q0�xθ�����f�bB��2X�^��V��g���S�0�*��� ��S���i�}�7)��5���]���������a�dOçbҞ�����Q
�s쨟g?�^��R�w��ca��T��)�kC�BF> Q�w�m'S1���=�w�߶Rڇɽ�y�X al��F�ն }2p�@��|j+��"�I�w��x�l̄�S��7��@\ם9��ҷcE°��܅6�;:����*3�V���!4�qÜS�yN���[�ϻ������a�G��f�ל��W�o����y�{E�DBɟx.|�{\^�cJq�o�@@�	�m��e|ijjx8�Nx�l}��@��S���X	�A�`��O94�z
@�;�nfN���L?f�-��a�5�(���H�U 3����L��T��/@�e�J<�pK���E�eutg @Od��R߫�^��/��x�.tp�f��v�)�^�&�u'>L4v�	X�(72J� ���z580(@2G�cq���#It� �`BTQ�����l=�� �#�sq�IMq]�����1���6i&||l+@4 :�3~��E�yp-�8��0a��h�������02����x���xBE�v��G�qq@�P6�׋���)�e�.�x��ʹ�V�#�ZY8�Z���l�pdB���t��`�!������*z:ʍh�y��Z���o�Qϝ7W��k��ФC�F5��. Q���3Rmkp������܇��r9�jˣ�Q�6����1�u�����b,�%�sB��©�S� �%Xd�
�����f*ӳN�_m�Y�P� L`�/Vl4���h�6�P�דAրɛ�A2A�O�N�Q �6GwC�l?t�V"P�d�r�^�,�a�&��<u�����[}�5NF9f���r�����] 0�߾1� @�@�Ą9�}��	��K��޾s���W��W��qJ���	�DT5~�;D@�68?�9��c �$ ��$>s�4�#L�;^}E]��2J8���MV��mSWm��(~��������?�֭]G`��'t7A%4�+W���e\@l��d<+$�^���$��t>����ѣǌ[=���Μ>�~�����͟�n��f�?0DG���>�,A6Ώ��� ���	mT���a��@�Q�wh8�~��2��h1 Sٶ�	 &�FPd�e"8��	���F��Bp ���cA�N��@,�k4Ø7�0�1����Gl;��Dh����MUv<�m����g��u���N��k$( ���o��Ll���Lk�,��e��'���J�!�q��
 Ӟd&%}1NA��.�K;2j��������}M�ע�ʯ�h�!���'�wĀ����hzg���_�C�ڙ�*2�G�!#�.Z�
�Tf�y\�-�K
�ǌyat}e8�`ɌP��I;Q�zJr͞㇠6�St2^�����2�G75��fVUk�)��7��MU]�Qw�}������>p����,��-����h��w�ܡ~򓟨O��ԭ�E����!� �����`ZG ���<��Cu��q���|����o�J��Z�����̓��7Z��x�]L!@�G�����wP_��i;v�������� a���#����G���h �����.~룿E?d�5L�Xa�I���2�9
��8�	��~������"�ΕM@(����b.?�Ѫ
.��7<�A��������,j��oi�5��,(ь��m�\�V\�eYs�,��1�i�#Kc!�gc���2��"3R �熺��"�9
n���'2���@�Pon^�
�J�L��Nv�S�l�(^+��n\My��ཤ���8|�9g��N,v���	�^&2��J:d�X[�U��Zݬq,��c�	����S/�(8@�f�|!�Cd����I̮�]��{�����
Fk=��X�0=oy�>�����n��Z���^���-,�`<���T�Ώ��D�)>_�����CID�[��۔�޵�`�&�БA��;����l����QC�_ n��g����R�t5k�L���č���9Ca�M`+>����E6.ji�/�ò���]_߃'���O �̮���x'wL���nR�Y5PSUr���ʪF���U���s͍�L
�Eo/s�L�|��/�\[*�ٶb.G��L&�i���];��EՌ�TOo��ӧԑ#�ԕWn����#X�3g���N����|�(��+�_�[<pT�R�U�x.�ׯg6z���Q�c�<y��pkk��f�f��O�g�}���k{v��P��5��׬��A3�I��G���s�n��@�v���˖
p~\�����$H\1k�,�G��������HhVw��u�С��_<E�,
 �GFr�f�9y����������Ѱ���um&^��Wjh+��+�G%H�죎��wtۋ���>dLR���������e_$�-�뗅LZ�r�0�
���iW��l�@�['N�a߁�{\��e�?����M ��m x�˸�]q�P3O6ז/��|~ܔ��#*�H��QYW��D��#���S�l f"Y�����4(V~���}���gB��=�B����dv��cV�� f�z�}��xNrMY�2p��k�<o9,�������!͂�L�XA˶��1�36�c;�1�fW%!�e~���,�%��3\�j`x@5%��>]���ȳ.0��-�lK�y}ɲ�~�H�<����W$=U��2x/��U&�ZZZ����a�dZ�EެGm�
�li|N�R�z��װ$4h7Q�v��-+�0�$�>�A�(�v�5�
d<����l����5�F��땣�/R�*�je!�%�O*�V���0ث円UUKV&{GG�#�)Mz}���q
`,�e"3qf;v��Q�`(�l�ӪlP}���'�	K�_��LJq��F��`u׮��I 0Iz�ujh|�^Sk[��ۿ�[��/~�@��a`x��()���m�ݮv�ޭ^|���N��A�[L��!� y�Ū��� �r�cǎ�y�a��/Y���@���n&8�9�̙C��o��`���G�,> X���l&X�O}�Sd�,�{�	4�l9ڶ.T�w����ཱིml^�����Nq���n��K�p� `o�&KV�7�*��zGr��s��6+��ݨl̦0~#N�֯�Th5ſ)��M��ؑ�G0i��j1���7B�9�͗�I.�v�g�P&2���?`wY��G�x��~4�� �ҟ����o�%��}�)�{��me�;�5��x��Ԣ_���~ڃ�����ь��Q��y�Aq7dju��(��}�y�R�b1vy�C`T���H�0��H,�{�(���,����0����sà� �5�:��yQ�� �mH>6uيU&W��?����To�G%a�&�����fA:R�G,p������G ��OV�2� mU�u���&.���F���}*���|A�8 CN  ����G��� фz�՗����k�٬������ꧤ u?g�28H�q��>�X��F�H���w�n��պ��;�>H���z]yf�*��0����N��lL����R̜���k������;�x��Ծ����Ԝ��ղe��c��d����u��g
�	Bb�g��q7y�b�(��/�^�XVvP2c����Lo�2�.�d�J�����nB;Q���*�\d �0aQK�|FLduV'"�>>��C :��0�DBT���Yz��<���l`�|#d��,�H����ڋU�X~�HB<_/�m����F�����L�ΓTL�tL`�O�Е�уS"W�Z��������j��@���L�K�Ȋs����[�Ȭ���k�5��	���Mϲ�vSft�����h�G�� �2��^% ��E"
�Y8�@�Q�'0q.��P� ��|n�T���P�D�ȸ����&O`����4p8{ꌀ[W���|_�-�TB{Ђ�JOȲ��)V���v:����o�/N�1��E�Һ͎�6�'@�?�)^WgA
���7~:�:�� ��d�p]HF������VHK�{�� ,�B�8n�I��������Q.��_�qK5�AR �vȹp\�34�`�!Y������:t��Z�b���;x�������y��/T���w�����-��"�z7=��~p�mm���z�z5�kv�_�l�5M��J��b!���NVl���I�sQ�8��W���-����+�?�@Y��SR�$0��"짲�j\ �/��������v�^�#������F���n��>s�.�=/����]�XH2�~�)������E��/�:=v�Ւ.+�]�.y�_p\gX;���1��55�_�ཤ��_&�Wd�����l\�Y�l�Z���e"pK��)?R�3��X���5!��*7�Py��D�=St9�-s_k�08�r��1q>���,=ccq3ɜ��_#>]�Ga[��XЮ��S�zAI{�&j�x\B�<��K^i<�oX�<b�{����� �a����W<V��|����$b�BQ� �V�`% �A�
p�z�=�]V_��n�`~�%����N�NO�څ� ����:c�_炪�GƷ��1�C�޳�~�YZ\Y� �JfOC���U3Ш��SZF)��ʁ6S�	?�.�q�k�j�
^��]{TSse  �����h�&K��R���:A��9s���_Q}�zԉc�����LV��1�:�E��>���.��'�xB�	��+XY\bs�4J D�׆�[��@b��J_ึ���p P�+��H*]��?�,��_�E��˗ԝw���QH8�����j��ݔA���űaIf�\\��֭_�ҩ*�]�A'�pnt�8C��+ s�<���5�lw�6H�ݥYW�`�W�I��N6�1�!B��W�zL0��v�JM�3�F�Pg9����Ym�U%m�p��򙄀�q/�N�[Po\�F�]���n׉Mp�#G�pG ����1�3����M�6���u�ܰ�C�j��ڬn=��[%x�ݥ�������v˟��>�wxca����ʡ`�V�v�a[g��<'�#���t�".!�ؒ�S��n��-jٌ���{�~���n�R��Y�<���R��ĂQ�Q4	9�+�$/�L��3x6�m�d���:_�X��cwH�H]�P(�9�!(ǵ�m<{��h��I�癊���E͙=��r���}��X�L��^� �%W�&ʪ7��1�~ wb�u��ꛙ�����&+z%��h���F���콓`h�{�l:���e����/�TVQ�4���=y�I`� �u�I�F�[S�B�n�H�DS�A��)�Q��x "ϝ�.���t� znR5NkV����/r"B���`����uLZ��=qqc����c��u�W�d�ܤ�2��z�ŗTWv��0�m�m��>���[���S �a�}�Y�g����=#�0Xԭ[��lru���L�q|h~����յ[���z���6{v^
,&䚡��cC���� ��9�k"!��G>�a��c[�?��?�Z:::������/�����Ƶ�vۭ<��e���S/��<e���ﱎ�|�@�3w.�`�i��`�lߌ��B���?/�M�vc\ ���~ӵ�wƎ�f���K�5X�Y���n=���EL}S��L����{yĤ�6��:��}oc^�;1�n*�Q��O�ʏ��jj- w��v��<�dA��B�$��6��1�!��m���x�<;&�0AÐ,!a�:��Kz��3&�=�Nؓ�w�s�e├��W� �%V��_���%K^��V�\�I&c�n�ޚ�ylě-�8Bw�!(��k��*:x���xbV�r N�p��s_H��k�u�Ʉ�����=c��F1_(�0jt4�=Ʉc=H]Mǒ�v\%�+G\3��nu��ᖃP�� �q,F��w�l��ݳW>rD͜ե=+�\�0@N��T�U��Fư��"����}&�}z�g��Ŝ����nuMj�ƫȜ��ԪO}�3�A�_cC�Z����[Շ>x]Μ:�f͜I ����T��-Pg��R΀Iz�L���y�ݪ�������l�Z����|�BM,�3���r���N�xb�
��ŋ�3]���`�r�&�g�0B0�)��q?��{(�@�50�8ߺ�kմ�i:k�\���*Q%�~㦍jQ�B�h=r� ���/ǰ.*�-��5��Ӌ��(�x�y��h�X*4��k���iv*�/�Y{�>�{Z�sca{�(���,P(�*��XR�c�����z���728���x̑�M��3if߾��Ǐ��ɂ�,����� �a���O��X[C��&��6��ٚ݇ 8|+A��A[����o��	�=�`��Z�_�x&K�شr�h�kDI?���&�P��kB���9
�`�	�:g��Ν{P@xg
�_���
,� xa�_WWwB	׃�� rm�/�M�4d8���^�:^װ����hq�;�߹��Uy����ۓ�MZl���S2�l\��z�D�l�0"�:�Ϡ������2�2i��/�����X�DR�ڈ�ΊN�� %ns�5�5��P�b�2��+����8�O�1��=�WAA*=�w|ð����x�F���v��xc5���̙�N�>M`�����F������ ���dK-��"�Vl_�Jcj��y��V�����Y�p	��:P@�P
<u���pQ����9�	e��.$�\�;X"X�Ἰ0������1����%Ƶ q�,��ܹ���� .�<�����W�TGP������ů��~`����J��[ޠ��F>�w��(�Y�f�[���8Ƽ�k��/V��㑧���p��3/>��Q���o/����&��q�QY�%��MNx�͌�+Q�k���WŲ��g�̍cT4!�-�e���T�P�?�J�Z���G�d���"��sb<C9Q�ef'~_�i�~���;����4��&#e)���}���-_������i���X����&��YX����}{�@̔ϏQ��8zp �g3=$ʚUZ�`��_�[ƞ7B����+����NkL��!������eYo�<h^%[.�^\��K`���Y���|>w�V�e%P0 Y
��0�0��������_�+Hx 'S�б�7:!q@7z8ט�CUg�t�D"��������p�}wKF��LQhg�Aw"K]�G�eMʯsK�V^�ي���&�g{φ9��PW Q`+p,kق�֥����1lΗ��R� �>Z��[@9��TBMkmQ�t���0<
25r�OM_8_�z�L�9
P�t\ Cf<�k�m�@{�\^�w#5�������5���V����gmm6^��Ւ�DI] j�V&5����EE����F�3�vP��rRo�|�R	��a�N���!\`�EO����5���ur��=}x��>�ٶ4�'ذ��x����
</����i�kQړ��4t�E�5*7:�]�1ioյYNй�0���S'#�Z���g�c��s9|� ��+��/���C� ���U�/_���m��˗�����u�^݂s�t��u�M#F�+��p�> �v+�� @��ݦC�^�t��l�?\�E�<54�ڪ������h铃�cf��E�#�ec���8�G�q"�L�ﾺ}�r��jl�!;\ĂSƜ�q����l�c��\Ӈ�xcƝ��,�
f�AY���>[ʗ����Z%��3X4}R3� Z£�Z��?9�O�mִc
eX�ٱ�5��=օ&�+�k6��������EQL�b� [G�sї6!�"S��ko���JH0�T:���PW8q��[���>�J�ƻN�w�:�����JG�*Y�m�Đce��M@jU�A�И3�C��Hk�6��_�j���	�כ�e���e
�^�ł�d2���=��5Uh���8��ݒä�#����ߘ�l*NmI��9!�}s����+L
� 	0z���5���F�b흰ɕ^��~W�ɶ��J�m�MJP3����AA�to�ح>�yk�p,�`I3��6
�v����+K��\�b�\	xY��~^?v�ཡ�^�ƔP3"�[�Y?�Y{���0�g� ��	��k6��Z�*0��ēXk2���u���a^v4�p P&V��y?I��X�R<o��g�Էk�.2�V���T���� uf�ύ�	�Fs9Ԇ�&��pN;O� �o�MŢ��)&�o����Y�@H'�� �a_C��H�~p S ��;^���z��{mlhP�C�ղ8}�45�`�?�������}\/���O}0c$Ӏ�ٝwݩ�?@��]ǟ?��F�Օ�61���9c�t^$% ��f �ƍWr�0�?��e��	Po���I�A���_���|��*+��E��$�4���e[���oT(�)i���� b�א,�d�(�kq�2�	��.�d3����^�c��F���'�/��9�ˎ��K�C�g���̘�n�`ȖJ���&Ṙ�:ev�,S���ŏ�G͂N.�@��q/LuɈ���,��Jql�#4)y,a�_N�Q�>�Ťhi���N(f����簿�\��\sS��t�1�oS����L�K��o2X�r�456^=88��8�c��2�c����d��*`�6
1���M���U��l����x��-�&O[s����N�q�x��i�����w5#��Cq�}P���'���n��d#�	�V&7�Kp����:�1�c���cs}�O���K_�DKװ�o�ZM�I@.AZ-�o@} č�ˢ̸�o�8Rn`Xi��3$p���=���
�F�A�B�]��9S��O&��
d�Q#������F��Xq���ݴ|�e2�a[�
݈ �a\/��j�R�i���K WU]%@�Agƒ9�L�i�����u��ij���<����iM����zf*C9y�8�? P�`�w�ܩ���r�u���nԱcGB�3�\���tR@]#�"���2���w]}����Ӫ`�R�XP���\^;#�;'��1e�e˗��+Vp��w4?���:�����X;4>�� �����m�-[�����x �����wߥ^?rD����j޼�*'`��n�|A#^p>\,R~�-��/ @a���Ծ����@]"H6y �]v���:y��, ��`?��t.��`�|:MKyU��:o�e�������a�<y�h7K���� �bkG����c��>��M��3�����O�3&F���G����� ��&�곒(r[���0��X��ԣ�����t�4��Q�-7���N�*뒱��r�$�$�:�k(+v���c�1ڮδiҨ{� t����h�5hw��%�˕��M�W��VY?\�K����*mܴ�2���r�)�{�tfh8�)�������ŋ��H�Y��h��NL��O�@�(�2"���r� 5��lf���,��e���[������i @Zn��zGE�+�1S�I}�5�Y���e��S�6�:�ހ�Lvr&�-ÅX2��0y�I$Z�x��5�+��[�8�ظ�:|��fQ�p*乍��6����j��.U<������A�m�V�SRi` �v²nQ_+ ��W�d��C0 #3f���D}Ζs<��㪭�U-X�P=�����p�{�ܺ�����b"�l��x>��3�7W]u}y�[Z[�֭��w۪HJq�՚�ר_|�>���t��Vu��7��ә�/�f��4�h��m�6^;�����o��ھ}���c��ׇc}�w~�����&�.tːS�t�&�6 sڡCG��s @�7
�7$�@0�l���z��k�๮^����<`��b���9Lַ���Vhg8���+!�+�����# =��租z:��T����z{��|��q�k�NK��c?�^�([OS3g�`�#RO:R�@�ޚwm��@��a����Kk0�{f[ZЎ��zƎ�$ٔ��8�d:U�&=ioC��F0�>Pe�Y�%��Y����W���zb{���1��#C�L�$��k�1���������O�q��:N�jw,��#N-.vM윤�^(� ë|�T%п+��p�����4����(?�q�IqA�k�6�Y��������\�3���i���r	�)�{I�r6��`�뻯�f�1�d�q�׫�Y�}����  �$e1�诬V6T���O��&�!*w�^@ 0m��$���	貥`l�pL:\�G��lr\��M�qXԧ��QZ����f��щ>����v+{���m�����\�P�s��W���*���dX�l� ��4Y\3#�U��4�,�e��?�>�o�����p�$od\���J��p06 =�k��mx��X\����`��1�s �9�}Fܿ�ײٌJ;q/���q���l\���*������>��� o,��U�9�d�g�̀~i½��%/�ѣ��#_��z�I��{>�Au��j���kT__�� �=���==gX�S�7]��=�vlY}�[�Pmm�v7�j��S�(� ��׮��F���V��P�fu�-�`�"Z��� �`����z�Mj�ƍ����:�ӭV�\�N�<!?�$��z��#�W�9ӭ�z�Iu��!UW�r���l�?��������ٻ��+V�P8D������kj��ޞ�z�J��;Td��
�ܿ��z�˖]����G�غU�C�"s|,'����ݥ�,lr*�NP��:�S��9��r�� ����vra1::�F�p��p�:���r}Ө����U��l�ԏ���JZ�>w�l�G~D�ٽKmذ^���w,�4i�^t�@W����I�9��p?�^?ĔֈI�ɔ�
h�BZa`_'�˫2Y�;&aу>�@A*��r�?0q 6&@����I؀�2�[��X<�S6��,��!�/�U�?U�6G�G���2Lg�E@N�����JX�x��C j��h����T��MBt!f�L��F�X�o���iYe=N��8e����d4M_y���gv��<���� ��Xø�3����	�.f������8Bx\ġMC�;v��:��֮]���B�[?O�s�8�nS �}S� �%V8P(4	�J2��ͬY�_>~�X,��h��ٺ�V��XeW&j�Ή����/Z*A��&_�S2 �js';�9�k�^�n�=��4_�o�Y��
�]ʣҊ��<�+��Q�Чb�v�wg�������N������6#7�'s&���3u�}��v.T4���9 �ˣ��	�,~���dM�4xV�ܸ������- �!U-m�QC�P�S�D�X��@=�G�TFE"�v��p��RW
0x�x�d���L��j����^�EF���o�o���:u� �9|}���W�ݧPx�h����VK�,� `� ��,nk�\��/[�dC�Cj׮]j�����������bZ�2� ����;�;�,�2��O
㪭��SU__K�����ȁ�~���5���xH* �Ж���r��1^�ËkF�X���q�EA)<���l	.���y�42ǰo�����>�jdq-1v't]H�9s���D�8���q������pNآ!�.-�u�<0Ы�Uib(�kNɂ๣�Mu͚!`Kk��3��ꅷ��{dR��k��{����8��#�,������}ft5!�y��}��_�����N�"��|�� ��jx�a� w�&qM�X��^�N�?n�*m<�-61�B �����t=��8.&�1u�6����J%P���qc�ݭ�,��Xr#�&k��P�m�<�;o�B����~YBR��փ�'��X�r�V����T�ڿ�2x/�b�b�*C�7,^����V����ӧ:��H���r���ރ2��A�Z� �<d�p�G��`G�0�ۋv��5���>n�t�+ T^�D�4Ʉ��X���>�Й��L6�Az�
�e]9��H_�?���J%�ÄC?��iy��m�^+���F�L+%3h@��6	�0d2��͟4��ֽ�����H����K�N{\G܀�	cb�'^C%ä��G��
d������D��O�~��~�Y��sL����:���̔:v䨚�t��i�
0)2�5�2�vL�b�T�. n@���Wc�a��)�B�
F޻��l���5o�u�\�,|\a}܊��$����{0Ķ<��j��Ι=G �N�$���$�u��G�k�Su�u���Sv<��C�{��)&�8* ,���s�� :`�t_ݵS�򪩥I�윩����g���nmk!K ���,u�=��ھ�%5sf�� ��լ�N�K���ٳg�ǟ|���v ��)FO?�cGgѢE� ���ײ�� �n�}����o����v' � ��5!� �Z@n:�b�9�g ���AطO5	؝&Ϻ_�/%c�B
gy�u�ĸ�dh���qJhO�l�ϐ8�Y�W0-�7F|�*�w�f�]A���k��p=�#�5M�˷}c&�J!��#��of�K����m�k��D��;&1�v���Ay7LEv��ZLE���(ZZ�GdX32鍛H��Z��q�[L���ж���AfW&2f���2�u:QKN�:ۥ�L�7HK�L)<ƹ�d�,I_���{�
+�$��W1���D�����KL�R4��8g��ʂq}�C *�}mШv
I3;�����������P(�/�u�QS�}\� �%X�,/���˖k��m�������2'<��,���0� &�-��hؕz,�_��%@�@{2y=W�<2x!�A�lܟ��@lgc� �����`�c��ף �u���$M' ]o�t��}`�(�� 9��LD�6ӫ�G��K��Igj&Sԕ5t��Ŵ���irɺ4(c���C�c=��(�;8`p�@�FT:���E ڨ���L�gϩRn\%eq/�sK
��eP�ug��R��КsZ9���h�}�Nu�7p���z@͚5[͘>K��I�k�n��#?5I⪽m:Ͱ�,J�~��X&�UW\�Q��S[��Bm���ނEYs�4�C�^��N�fw	��W���]����0��5�ZC�-�FH�ˍ��Cp[S�4DG�Ժ�e����זNWɤ[�r#��q�z�򗯨_|��.���K�|Y�߿���3���E����� �믿��n`Y�oU]��>��N��fǤ��ޮ�z�I�(�X�f��%�E���~�s�,oڸ���������O~�v�qq�&���靅BQE�p�m����؁yF��'����k�	n�Av�_��2���Sf��jGD�`T�$�C�0. ; �1!@B% P٦zU��[��c'���2n�:�-��y�!��`w�.�X}��U8����{6Ű�F�}'cB�$��خ��ʥ��.�Y�qm[YY�)��OK)]D�͘=S���������8���"��D��7A� ǐ?�;� :��ǳ�d�C�+�b0i�[8gJ�<4�O7�;��2��t\ƟZ�t�@����hͧ���L�K�7\7����+et��k���������7/�8�`��ے�Y2nQ�P�?�+5`2p pN����&&<�$��Ą
�#je���xF?�t���'�d<��2��k� t�6��9�e���(��p�h]������U�D��o�K�
2��蓋�4�6޺`��6�`Uҫs���&�| �l�,���^,fKP+J��`�dm�:���XtX?�f&|��k@&^��BOf3�����2�)w)��ڀ��@����F�D<�eu��Թƪ�/'�D�@""5���k�L�ͱ�f���N����j��՜ܫ��2�	lhoQW^}��ѷ�Y%�I�Q_���~P͘=C��9����.vt�5T�	N�f�%�֙� N�-[- �K�i+��]��fjv��մ����+�!	����7�C��J��l�� 3�m�r���vu�G>�~���������V���k�N�,��f��v�dttp[) `B�͍����}�Z�>�Μ>K�-�\O���{����{Us�tNЛ6_'�$+��Sm�x]"ɴ�ol�Aa�;�� '�AO|��!��\��R0�kV�&k��piT�>}��-Y���y 6P�<o�\��&ϭX�\-\�P�����e˨̈́�Ap�W���s��P�v�Qt�`@� 6h�?��?���`߻��;����rߺ]�ս�~8�i��9�%x��w�}\ �F駊뎹:�gKA������[�ZǛ�USZ ��~5&?UJ'Vp�����ԺekU�:�
���d�E�N�=��g����`}z�t2��=�;�Hgvz�����pqf��ɀ∌���2��ʤ��y�	F֠";S������dZ�:_3��j�2d����8_M}��7����l�d�k�tT�� �����*��S:�q�&�я~D}�[�R�?�x����=�g��s���d=���|��_[�?��W՗�����?^&i��n Y�{Ĝ����P3g�T_�ۯ�������,@�%D���?���M�	b2�;:d8@��$}�ը�����퍌��٠���!k"|������e����;n��-�ܲw޼9�}~�)�vS��[� �%Z�p4[:mڴ�k���y衇~  3�mTZ'�?0:`V��1I� =�c�������*��/ w`�z����/�ikm�m�"���T�`�K�[�ɂ�~��B1\e�|L�*�	׊A  �I�2�S}��Y�������c���k��3�P��	�����An"��?t�-y�� �� &և\�	����I�j�����`�G0�%�6�5�p����t&d\3�].�����z�G?V[6oQ��|nL&�QN��?�Z��'-c#�vzN�V��=��}��3�4��^ .t��N��ld��OSc���mVg2�)Uhj��jku���omI��V��0�}A�	�#1�F{��s�S]]��y�ͷRN0>^ ��g�%�I0qK^�[�A&B��`�ƶ�F(p�r�-����)my��N���sט����՗�g�>]����C���'����Q���%��lc�4��U�L)�p��{e�f��@ml�zbl��(Ԭ�#������� t�  ��V����:d,���j�ҸJ��"Q��nt�����|� L�ۮ�Y�s�'�ccc��{^�#��&�i�����"��,���A��Z#����匌2}�pO���|��=��zLg�t������5Og�& Ģ!#���;8�`�@2J��.�d�;&��z|솋шK�{]��g�<��C�M X楽Uɢl����˖���~J;u\��3b�u\.hq��c�sZ�h��җ���O�V|{���2$��؅} �g<��������տ��/|.'���c�Z�[λ^my��`��|�wy�]��3	�$p\�"{��5Mcb c�+����	v���w����g�,j:�v��sp����ѮV�,C��K]�\�}���fu�z}��E��rQ������*�e
�^���>V�b�O�`Æ?ٴi��?��C�bn�A�A&%�LlCC�H/X���vO�5ۋ�U�4��ƪF502���l�V��8#2Q�9�n�x��[��]�Lm��Y]S��;�B�Yh�d�IfA��2�p��ٯ��U5�) ��yڸ#U3�� O��qn'�}��c���ۓ6�2%d��sP�i2R�G�w�G�<��	8M �Y�, p&���&�ly�ve�l���h\2�ɭ�t2	m��#A�=�ec_4XG[�	d_xn5���)k�Ke�TUC�,NF� �s'N�]��
��())�}�s<˦�[�Ɲ�t҉��h�����)�wuZ�r��^�Ȅ><�5wm�m�p�'m�8h ���9Ƕ���F�v0�VsAW���U�VQRP' j���U�6)N�}
���>sΤx�u
X��c�Z�}=�MkU}=���\TUe,�QεwTp�[�\'mLg���:��Gr9���z�s4��I�-N�g[��>�~���1h���N7�E0
�Z�C�2M�.�`['�˲����Ǘi�çl|\K:�8`�[�B���m;k���| -�3���ק͘A���
����p��E[�b�H��E�=#*8J4����I=�3RO�d�Ki�n�Ǹ8�1XBY�������A�]$�[���ə���+5���=���x�Y�MP1\.�:M�_��xK�-�����}��괴��7��ݸT��$,^6n��-_�j���׭��閛������͹���3�>�T7Ȣ
�z���>�῔�ñ�w~�/����W�{�cH�U;2 M6�o�A�_0�;;��ڤ�|�Iu������ףm��AɌ���c ���[o������U��[��*�A�6�y��C�� ��,��Ӧ5=&`6'��۠_+C��é0N+S��]� �%\8�::;U~�Qյ��-������g�����g�P���2�9 8�<�c�� ����HԚI<NiA���ۨ�/����][��ך�cp�c�1$5H�
[�I�@��|�rֶ2>'El`�� Y� x��`��%jߥ��u�C� 	LpnIG>[�J����iƬ���:\�O���B�kG�[l��� m ��8�7]�f����}_�h���f����sT�`>l�3JX3�LTJ`����W����٧�Q�-^B����`��v̝������½#Vߩn��˨XQKM��O�8�]�o��~E0\2����;y���SE��e��q{�K&H�h�</��`Bfblg�IĦ7Gig`baO6L_�>�+�l��@���3R��Ϻ���io�zԬ���x)��cd��n"��6�q#m`�	�9Xl�E�n�#| /�P���gϒEݠ�e�P�#��v�ϓ�o��d ��c\�e� j +�}��Ӹ/��LL���}�#���+u��N��+׆��w4pNȤ�ΙO�/e� 0��\�y3�.ԗ,���v@��ܸ�K?O�"<?6�|A`z���  9+`�Ё��ˏ��k5��L�ZڎC}8�V�-��=�9��5cx�?ܩr��ۅ)'�)�]'51h�,�Q�d~�2�o���M����-Z�h���>�bŊ�ݻw�h;�T.h� �A�+�6m��z��<}�Iy���.�~���G����{��I`�544�4�ag�k��[S�y�����A\�n���}����q"h�h3,T�ׯgvx�w$H�ks�9�.�4hK��l�XX͘>C}���TK{rp�w8۞����/ٮ06%�6؍;����H�߸�<J�����n_�3�6�v�7U޿e
�^��n�{/�(����[nQ]���?�����L0%��2����7��ʜ�]���j�e�x���5Cd���uf���sȐ�q�0 3���ub�M�	sfW'1f0J%tTy�Q5��A/���*�	(�,d�T?���d�0ia���*��"35��r�2a]�q#'����pn'�\fY�g� 5}��b�2��If��u�4��#��"5��r^�Q5�5������t� eq#�@0��d#��^����6�ky�-b��N��<��d\��fLr�ׅ��e�m����%���~�A/`` v�%�/�,B�~�_���Y;���p �/O�y����|QU5��t�:{���_���0;yF6ʁl��7����y˨���b!�W����T}C�Z?�b��:vLO�������������Y�=�� 7B��A~����_�F-�6~�X��_~�dЪ�tn�cD*��W���PVt���׭�iyI�
�1�\�# v��-j�yO�B��ڢO��`q8hҠz�(��ٸu���Y_���7��+C'��c[��իWSv�SWq�� �S�NL��gu� üm��6��a��}��G ��O��Z$��;t�	;p̘Y��|m��'y^�c�^{�,���h�(%SXtC����b�]mߥ8.5�p�q�.?�S.vf�.��5.�j�������9d<�@q�o�~��Ff�֖fS�z��T̫d,5�d!���zk���'	��`�&IPڽ�h�lc�s"�-���-�x�j���mZgN
}�� �l�N54M.^�²EK�oj��#�V/_�������g�}�WZ#m��j��n��������2��r����K�-��������տ��,������)�$[X�t�_Jz� ���~���/��O��ۅB1�<�'ߕ��_�~m���Ӈ�����6�{��:|�h������9&R:�vid~>��ύ/Z��W��c��#�,[�<s���Ǐ�B�i?qW[�z�-��U+Xo ����C/`��������n���) ��*S��/6�Ֆ�Z�r9�M�}��1���$�/�a[<���$��$�B�vC��˰�`� ��c�X:��5k�3O?cL�]U�+�h]  ;����}������3��a�	�pJ��Lp�a�t�U��W�HJ}�+_�3� m������a�C��5�]Kr��q/i���;�oB��:��z���j�ܹa6,��}�v���s� fAuu��l��~8H�F�DAp.� �r^��6c��@Y2̒FR㣉A��ɑ����&{���F�� ����*' g��W� 9j'�M	&V&�֮����Q����!�r^���bF��g �q���`��A�d��t&�F����Θ٦�vw�u}��s8|�u>�ٳ���z�3���jͪժ*�Q���ޠU�j欙���kG ,a���3��v�2l��%���	���6a���}��|��3gNg�=���f��b��$�q��Iu��ABH�]�3��a��*����ѧ7����7􉭭-��P����2��k���mhjd��� ?��*9��_�E�/_x��
��,��R.�ǃt������ѣ\�Ϟ��	�y��
Fy��_��ٝf�&3�k;}�e@�����7�-��=Cp�1���%#� ����#�>8^NG.��fsdq�s��|!������Xز��Y����xy�<�C��������VfyZ�\���)'x��7���Z�i�����,�UJkk�� �*L���s>���t#��'_��'���������\3^�;����융�;?�G\���Ֆr�gTI�J����
^����K��ݳ��?��Snb�?�tV�\�~�m?[�t�#H��`_�u�T¿馛������?|�<g'�+3�Z[[�\�|���:�b��	��Y�rŚ{��^���U{v����'FGs���U�V����w���џ�O^�A_�m�����SO�wY�M��!�(���s�^ǈaA�5|�u�&l:n[j��8hI\�K���L�߰��J1{:������詧���/ݺ{���ݻ�.g��*V�H
�p٢E곿��jÆ�/��/�_��r��2��
��P�|��^�n��md�~��V�sЏ��nA5�d	8�J����պ�Y�;����$������?r����V�q��8���I�}�tɛ�:�\{���&���,��s �&W{ ��$�����y��m���뽖���w4+,�8�3�d�������D̫������s�{=�-���zJ�	�)vB�F���ݽX�����E
��8�k���1	�����6J3L�����	�G�[,8 ZA%l���j�ڵ���D�>5y�GO�����mS1_k�Q�&h_��<d���^vB "�?�X"����ŋԣ?yTuu�pZ���~��Z�?�� V]1�ξ}{�gw�T�_;��|�)������cǎ�_m,'~�=�d�e��$��.:k֭#�N7��Py@�ܹ�7hX/_��������G������E RÛ�A:(>���@��7�Q�}�=�8���5��}'���`�n�A}���W_%�����v�����uWl`?��4yM���S����3$J��l�Ŗ2��?~�l�8��� �s�eK䞺���7�� ���� ]�݅���a���_x�c�Ρ@���yȌ��<��s�)�c�n��@c�\��ӣs�8u�����eF�,��V),5q���:K�~�yH�1k�LY��` j:��V����)y�H��%���d�t�{����\YxүV~C�����J[[�즰#ȝ���׭�z������cw��&�y�Lk{�7n����� pʁ������3F>������w��O�,6477g��\������\>:��?��j���*�`tG���/������?~��l&�yt�쮯m޼����6Y惴��8Z�������m��ǖ|�k��qi�����Fda���?��e�8-���n���1yS����o߱�տ�g|��&��nj��K
�9��IN��ŵKM�-��,5 ��h���QS��[� �%^�B1꣈��
d^ VT��^�U������򙿓	�ܲ���4�3d��V�u�]��%�Լ������#����!F���e&� `R�����q�jS�}�C��=C�LT��r��q3dd0���X�_�zU�s��7֥>����0�߿��������^�.��]�|����; ���@(f�J ^�����s`���'������^2u�c���_�Z%�>��|�	��"�'Tū����1�J$=nR?)��=ϫ`��M����}ӁV�I�����٭mV����&)�
�u�w!h�F�ɽ~����o����舴�8������kV�����*U��R���v��a�hV�fw��[d����(P�j<���w�z�	 ��1�?��?Q{��t�����u���ܡ^�/@/@3���;�����,<������Z�޵[m�v��h� 
�@
��^ۣf
�(<|�Z�b�����9!۹f��꥗^PO?�$�ɰ(�v��L��0�F�ՙ��
��(�>��\��8J�3�׫z{�rw��MM���p�>����ʉ/�<�.�|,Yj!e�����>�%`q!��h����e˵�_�w��G�+���(�V��]˗/о\��j�,4��m�����֭��^�}�+/���#�G�� AC��.�t�8.���]-׻� ئ������528�Z�I6�	A�(v|RҞz�@w����USM�,,���ר9�4:�	85����X�!��׈�K˘�{1/>�.c��T��u��2./`��X�;P�n�n��P�U��f_z�.d�z�6�ؕAb�������#�
��,6�f2�w�}�W/sHm}�:{��Vft�`�߼�J�z�B�+����'NT��x㍍��Ͼؗt�����$&�1��2tuu����?����ƽ{���M��*�{���ږR���I	�����}�e��;_z�y��[n9|�u��^���y��5I�$�ʕ+�H��G����x�#2�_�������mInvkZK�Ň^�pA�m���6�ڻARL�K�L�K�������4Q쪴��^{��j!�ojn�{2�����~008�����xf[[��}�CZ[���W�.Ȅ֣J
	�{������#I9�x���޾޸0%�y�Nd�/�����p���յ���X1sŕ�o z�SO=�VPa�۬5u���ظ���pf������U��>�U�����=wN�'>�����}��O7$�L�2�`��}r���&�n��n����?�B���^����D6�N�_j����/�lٓm��R��Թ�ޞ�����t�#��>7��|nl||�hn�]&��D<qN�歵5?u��	���s#c�L����eڦ����xnt��ɘS���(������0�'C���R�пX��Vfr���TR���7�Q�S6)V�x��S�lH � ���p���f�Qz�׏�/�Z�Uh�L~yD�K�{��m��沪�� ��S�XR%�u.��N�گ5��Q��{@��j��`rjഊ7���}^�SY568,T�+@т����:�������\˽.�ʔ��Ȓ	rX���u��y�Q �g ����'���@: ���e����<caR(��j���dɷ��A@�N�����C}�������QC�����l��9s�\�v��aR��آj�jT����ܸjmj%pS�p�"}tx��@�_�X�͛3W�X�L=���d��Z� sL���t��s�L��1}�ڿo?m������sa	� �1�P0�`�)g�v1*�B�D<��p�HI@k��}^ڒ��H����[����n�E�c��T��w���T��5����Ȋ�޽�|L�W['�o����`�����B���`�H=�
��Y�qu��)\.Ϡ.#࿏�\ ��<�D)P	���mLk�<�F���[TU{�p yʨ>�U@�V�����gϞ�Ԛ�+YwL��݉ �FYN�,4���ϻ���`5��k���i#�~S0�W@J <v�&���ɜ7/y�b�9N; �5u��}A܃+wO�-�mS㴭�iI����a���O}��Y�Y@㜩�Qr{������a���>"i7�+׬����R���^�=EY�rZ�A�(g���i�_����q#fdt1:�ú�A�6۲�����z,�=66ڍ�f,f��0u���"����Pr]ו�y�ru�4	�)�$1(�EK�x$y� 簜4�{�o�'˞Y���m�Hr%˒H�bI0' $�DFt���{��s�}U]� � �V�FwU�p�}��{�>{o�>���d)��+��|���jmo (�q�2����J�ޱ�������#�2;��W��~��7=5վ{Ϟ_�⇧̓P�:N���w��o��7�|�]�t��r�2����ի�_��_r���/�D6�É�C�?�F֮���;��Ї�X"�`��+w��~���܉'�G����ե�����Vzzz^��L}�?Qغm��Ϛ �@ �QF��7�|�g�����f&g���H$��K/�<{���f���d\˳�3~B
΢v�\vy�o�����L�t�`6��<���67n�(��X�
������bK[�R����m�vvn.���q��M^WWW�L&��*�:����������'>���f�1d� 2D�	29 I� ��hb)��Ѷ���8�XQ㼕�Q�gڢj�z���ዜ��$,U�{���44�x�Ȩ#k�{������Aưxf�(��BG�F��-���g��LP}�e�B�HV���+h4�``F6�G|OdW�E��7��󘂚1N2`±b�4de�����Ud3�� �T�����d��\i���K�h_P����/EZbm)�4mڴ�v?�<=��1q)�,��ц�������K/�D���Ȱdn�ю�Cbr"Ҁi�G�������{�d�q.Fuc�ׯ��<�سg�T����x���Z�������y��� 4L�ǁv���
�m3::.����d�I�נl�"S�p�?�����%�|��\�R�Wi�E�y���hO�H�00^�f-��瀀���	���Z{<MO���B�9�,��;�}�ګ��"�Oܥ��qɄMh8.���o�n�Ed�(ƬRY�\��`�*�9�j�ք�� �������1`w1pf��0������ģ��!�X���D����@Q�p�Cf^��-<Y%�I�[Z��2�gJ�_%�\:ּs�_Tr�
�I�DE.�z.���&�3+0���J)�w�
�]�!���x�{]�B���.�J�-��S#�\4 �h���',x�W_}M����Ͽ��o�����N&�����o��mo���7��jwwO^V�#�2K���)_,��ڵk�-f�����ⷼE26%8A�,�f߹\)�h��������޻gndd����Z���馛o��-��=Y��0��@�X�~ ���/?P�G���C��u��~��p��1T�p�E;� �������7m��U�0�
5�~�d�.�߃�l����,��1��m����̀q�&7U��^��~�Wxp�m�Xl���R�:$~��B�u�^%Ov��=��)(À.� ��|��\5U]^���wܤt=����$}�_�L���k�s|�e�
��D$J2�{~�c�����k/������s5M���ѣh"&�c���b�\+.k*���^z��i���� ������d1��?�}���4�@���?JW^q5��/"b��-�u�v�c��5k�ɀ������(V���GyD8� �}}��1�"k�L%h��O��}0�ɪI�_h�<Q$�C_B_@J���j��Ā������y�9�y�Y��Ce y�B�OL��z�)�.>ǰ�qz�m�6`EQ%l�Zq��.2$�@�E>o�t@��{��K/��m�u�6n�&�e�����w���ӈ�[��<��}�G� �\�k
0��v\$�mh{T��~����M��D���g�
���67� O��x�q+BN�B��y�J����R7|,��h`�y�jv����h�WO��쒧&�٧���
�w�]�'G��ŝ�K�3�ت���]�Z�Lc9�+���2^x7q����
x�4��y[/�W'�JQD�,�W��Y���a��������L��|�js,�=�b��↦K�i>���|�~n{-��=�����<1oW3L��F,��&v��}ێm���U�����[�\��zSn$2�v͚
����a�I�\Ai4��/�<]u���'G U�aKF1K�lFq簄���n����6xQ ��z��iJ5��l�b�0'���+��,2X�H58���>?ԱTk2�`/0~/� ���B��]�(�_<�GU��΅�e,��̔�ʌ�
qmCU�S4`�Y�O�?�{��p#�>V@�R�W�*1K�m#���ϖ.���~";(�j��v��x�< �0H�H&L���Oн��mo��YJ��11C,�:m��zj�A���ci.G'��m�̏��"
�ж.k�3@��r��^��e������c(l �k��О8.\O�+�k���=��Ȍ�Od ��j�}�d�1p���Z��K/ 	E�;vL�f&���j)o��-�eŵ��2((���}ģ�<*��k��Z ,>9>p�q@��>{�u�	�m�	�m��&�\��+��B 7���>�;�6/���x�ܹ3�G��ۆޮp����6X�x�8~8b2��w�S\�@; �w#���>�s43�tk�:�D-�X+m���I�x�;��|̗]vY�//���k�c�⊫D����
3j�.i���ȵ9<SO�q:��>��yj��U�eQ��W�d)�\�q�
my
`ut����?��)PoW�L��I&����g�V�V��^OԂ]��_��D	~d�ZZ[�XY��]�Xx��1�[e���[����v��F9�w|����YY� ŝ���>\.,��ȳ��#�;�"!��Z�Я0(ϗ��4��lZ�X�?�� �?"�@��p3�8�ƀ o��S����)cS =�Z�X���-22p(�SVܐ5غc�*�л,�}��cb]�\�>cwW;�ͪ$ ֭����ӀߞC|  ��IDATk��f�J|?��h4�c���ۙ��Q�[<ȡ�Ɖ(�+�R�h��VQp���R8�#�xF�d���%�>h��hT2hx��� �A|S���OT
d�߉�e�JY��Ƀ:��R���������ſg��V~ߕA`����H����w����sZ��h&�kQI"Y���uì-��%@�?�|�Z�o��kVXe;�'�/P ����I��h3��R���o�@-�_��W�R
d<q:��e�\�O���xf�|�$����9=��O� жl�F}}}���,���~���J(i������D�88�믻^������k���� ����!�ղ\����rh?n#��x���
;��e���26��[n�/&�la83���o}�2z�b�s�3b�z޺�455-� ; �o���.�\���w2@�5���/C� ߁�ƇV0
�p�����xrxX2�8��!�Wl�7D�AG��hG�Db"gl��(!�%���֭�}����������DN�y�^����Lw��`� AL&��%���[@#�11��eB�,8�5&��c�='t��p2�S|����-�s=̀�(��@�k���ԳyM�1�P��BV��(	���fEEy��i5�!����N0��7�y{�[����O�C��ÆP��Ԡ*�Y���BEl�>��w�4Q��F����Aqy]W��݈Z�������9׉��f��x�B��$`�y;Y��d�	��n_�qk�`����zs���j�͕�9���m������shE�i��9�
]6�ԓz���Jh A���p����m��� �o� �1�@e�U����$3�cEq����$�J����
 ����EᡄeJh�V<U��JhQd�*S�7x��.h���r*2�j U�C�x ��C"�x�fy)`��@���~%���2��L�j=]p��� ��c�UQ���H&������>ji����!f2��E*�aGG�σ��b.�>~������Gx�Q|O�Ț�d�B�Mr�N�۰��;��dl����\��2��Env E8Rd���d���T>f,ÿ��^�hXJe6��Z���&i͖�4{b���g�56I�_|�.�蠮d�R�2��T��UV̖/�`|ժ%O�3�b���=�M�m��\g���!�� �8O�b��% ��hg�A5�5��d��%+���E�!,Sc"��H�V" \cb��'�d m]�=������T�q���ذa�pu͵�v=��ǈ�V����@0 7��gl��ۄ��� ���$+`�x� sn��b�)2]�ج?[����՜6�BF�|���}bU|'d��+����]іӳ3����о)�R��d�bV,�1��Pp�E`�� mv*K_:HE�!�@#��l%��d^�9!XR Ƿo�+�Gw\p>Mp?	Ċ�Ey��w8��̠]>곻��[gA��Ȣ���o"�E\d@ٲ���>����e��(�D;Q @��d��q����Ǎ�6)5	����F4�T�xDc���q�B�!M[<Pj!��/����Vuv��Yؗ�Pvˀ0[���M$���@DE8V�=ϒ�_ɲ����X���G�΢x\��[�j���ΐ�5ڐ�">'��|�xP�S	��U�����m�Rz� �h������F��]-�W0#��-���'��.�p��[����X"�QnG�{}�s`X����s���0�[�^��F����x�Q�� ?`�*2��7���7�w>�{�y��-��ME�'7����6����#�̀����t��U�}�f*��g\�}J'��;'*Y]\�2���6�C�K�Pn E��ɗ�!{�A�τ6Ep��P�*��q)p5ֻ � ��X_q��BS���Cu��@.Nʶ�"* ��x%Д���i��2�h*7Q:�d�7-�q�A���2`@���4�^���OP&���HsL�Ne� 
ʉ�q��1��4�{WSC��� [�k�ͤ�4C���uv���K���z!� \�k���E)�i�\*�\6/m�>n2�>o�����/�2���0�4�����@X,��2$�l��0�n��N8�'ʎOҞ'��(o�#�B.d��c��R���er��T�K�S�j�Z�����{���nQJ��偧Z�e"�I�\:3Bmv7�Ƀ�����d��be)s�q�ɾ���6=(����L�,�0&T�id>�j �7]�j�F�M�$A�6� ��	�HT�b0[Nr1$����ݝ�E|-A���(D����Pap�<dyd��0�mIq	x��,��^�MI ڱ z�c�����RT^Ee1����vQ�#�h�+@q\�!�����#:C���0��ܕ�l�M�Yv.g�6�
��fyn�_O�ӷ��^;�S(�)�8��7N]�u�����/�YSs�F�̨8�4�A�DF(fG�9�o�}�=���}Ltb�FF��
?�6Q�yk�w��;4J�2ۓiz��z�g�}U/5w�)떅g�v2Ș:xP&G(����7n��[6S�8'2z��<� �/8�,��nRx��>�� Kp}�Z[d_��"�A?� ^@��2���E߁f,��࡯]���n�BO>�����1�ӭ��*�Q�K� nH��DaR��>]��t�5����^_ ��_xхRT)��|�=��n�����U�����=N����|�۷o��?��t��!� lڼ���������e��ݵk�J������O=���[��h�͛���c����c�*"nmܦ��G����]�
��W�@�/���MD${n�
�Ⱥ��0�0��2����j�]�܉Rn|�L��|~���?N�N����g@�-M�ΣD{�I��J5��1�'50Y��DFJ7��6:94,v��ςZ�J�U���Q���E@U׵���5&2��իBF_Y^���_aڤ�,���s�n��@��"F����}P����WY�F9�#�?�=pZ����#_Oh_���F4���&��r<�[$R��|� �t��!�0�SRY\���K�]�c�Z��K�{h��kY���."�\�-T����K�2�P�Y~�s?��Z4��� "=U���X�F"655�diVi���"�
 b�Y��q���
�gQ}�idwHIVa��E��|I7���́�G$��:�;�zzb���mY�!����U�M�7��r�?���FB��_��Xp����.�e���(�y±���� >���2�8�a�s� m �*rA�\�Kf��9��6V2^���?��������i��Ɉ�n.ǃ*��%１^}� ��;B-�f��a�:N��f�����:��d:As�s�~pbhP,kᎆB(7S��B�JтX��(���������.2e���7��$K��F�'�$�x C���Q;@ / +~7�yb|R�f� n�y���X�8�c?@��^C�wlb�������

�>D#'G隫�b�y�>�������bd��O�T��/ƾq|/�~A��
��ߡU�W��䔀W�����廄����M_��W�H�;�/|��&�q>_dj���&���Z-&��)�u��w�u�]*�Tɦ�plq<���� X5���/z��s�F+2�Ȭbb*��?�C�4�d�``͓74_�V�����q?�𵌔���Sp}��뢵�6S%����M�`�������J��O�e�_&}����=-�f]p'����j�Y+Z(��b/u�����P��eU�Pm�����2��{_�.�3�R����
_L��|):����Z�A�������Q	��;�ي�� ��PI�e��7��㼅w�X���x.�9� O�z|�ʩe�OW�f����p�WB�L��s4 o#���n�z�� Bz���fq��}�����!�/&���;L�r�@=Ա;)�Ӆ*k����lh	j�y5@�z���.i5�
�m�u�7���mY��O �����z��<�U�����������x
���B�9�[��{>
�|��CG��Gw��o��>��������Ռhz��Kw}����RT���ݏ=I�ݱ���2����4��$�$,�����+���������)�r�-�-�a<~��[�i۶m��y9��`�3=w������M���9^w�������-�P!�d����>Y]�c����м��/�cPB���l \ݶl�J�18�E�Q� �%�D���o����/�Ev�8^�&X��J#�a�����7 ����*Ǐ�0�a*��W_}�ڹ��d��0({v�y0P Pt�v�J7�e�М�2&Q/����+(�C�Bv��G}D <�	�h�h�c�.[�衝�<��������ГxR��($��(?6N��x��SI*Oe���E¡N��VSA
i�������$4�8O�^�	
�������P ���XV-�%=���>[[v�ﾦ:-��Ӟqt:��S-P��Z�Wr���3���LJ����CaZ��=��+��)�R�C�[$)ȗ�[���r�P����s�A�hďr4 o#k����Jgk��yH���W���:�4@Ft�"��&��U�B&�,4�|��"≎*i[/�I���,%�%b��㴭P����~�����2�-�K����Ax����L$/�b�� �5��l�*f{��Cp
B�B�Фkř,ki��oeP�H6K�KI-��Z��EY����'��g>)��L~V���H�ҪM��/�#Ͽ$�hn̕,����]��=7S��Qʉr;Zb�4CM�M2� �(���#G��T!W�'�|Z�^��BiM�R�`�O�!��dw��ukӒ@N���B��{��p;�0즛o��S:tX�q�(@h�r��N�.5��ŗ���ǩo�*�~���bU㕃���O=E������]r��/|��_i4���_��:��pNfI�ɧ��}À�pEÊ�����`[��v�m�ߟz�Iqт��� ߠX�)����C�H��RrtUk��_j�C��D�d@���%�+R��U�T��^x���r��x��8��R�ڷ�Gtw�l���zv���Gl��L��z����iE\�9�L-�)����Z�++N������C�c���yv���rnA��u^�o��1-�|�8����#��\l<?�,P�)甩��6t���ۈ74�KN��f2��U�̥-�i�B� rF}A�lE�%7d�@(�1�� �2^��ր����qɰ$����c��wz�,V��! ������g1=��\��
�;:Ë�2�1��'�����E��2����MY:�ٹ���������OP�v� KYX���:29NA���~�M���(?9K�l�|ţ�):4z�n�O��ةl�Z� �s929���A���#G˒��5�����������q<��b)d+�� ��VY?���0x� Dв��0$ɤ���y����!�"��?�[�I2�����g����.�] g���e�og��0�`u����
P����$C/d���{9�^�B���k�	���g�x.����O
�`�'ο�w�l0x�8'���}}Bw �^dvq-aK�X������Et�h��2��ϠO�������l�Q�0��q����a:��j�\����r��MǩyuMq�2T�`u��4 V���#�e�϶-��W���gK�I�f�P8Q9Q��5�޴_��b)aL���~Ţ<��ơ����PhО3af�P4N�� \�F4����c�4�ͩZ�õؾ����:�psu���X��R?��\v����
:���dU���1�P�L91�吏�L�Q��eN�x`~J{�5Niкt#�T/lm����b��]S�L>N��#72_�L�MVo;Y��`�����[�� (74Gl�=9>%5��b������-Wڅ,/,�P�~p��^pr����O������OӮ�gȅ
��b�H�d�z�:�;n�������n��NS���������
���*�3"U Ż��}Er�451E�6l�<_��=_��\N8��?ƒ.���^�����E�C�����ںe����-޼y+m<o��Rdp3ssԿj�PN�<ɀ�@h@�
͎�n�(���<7����c���(�A��v�'&$����O���ki`�:�g	P�Ç��كm�R����W�*�]����)C�<�K2��ɮXG�-���S�L,���K1!_��|���q E	�ԅ��_F��]ɹ��?@sA;e�=k�*Q��ŝU�i-LFQ���Og(�m��}�'{&G�H�R�l�M1�Z�������R<*f��
5;��"Gv�=ߠ���L�M&9�P�����N�s��D |bm�W�P�����p�qO����&��}�[�`��```�Y����JZK�ɽ�UL���@@�������!�2�e�w��p�hP�#�ۈ74r��_l�0��BI��` :�������ʒz~X����>5�<��\w����t����BQ�&x���[I����ڨT��B�=P����dzAߨx�4M{�:)�������z��L0����/��M���_�����mZ�j��
Ez��A�^����f&��k��]��G�}.C�8�Ю��]��wQߺ�425A9�D�HBL��OD�})D� �(@�YL�݌So�1�<����������=�%3jd�@-8r�(��Qe��@P9�y��^�ֳ�
X���l��E&�S�C�1�� ����p��02��;����f�8�f���	0��>��jKk��3@��E0�����`��ǵI
�@5?��O��^^2���w�y#������� �*|�b�Q�K��Yv�N'D�O�%1[�g$��p�1�����&�PWs+=u�wh���J���S,��i�.�I�6o��'?3A�U��σ@�+28�d,�>B���@/��R^&od0����yƀ�e�,D�[��֮F��84x�>M$n�9����W&�ZAC�L6ڪ�˶�%'4� ��x3E�6��eEj�.������Z����1E�jl�)��"5�ɭ[ �y�7/�[z���3v� ,�u���T2Ua��-�ƯY'͹�����4���V�āC��/���%�Q�d����{��3�&�N�(6)L\5g��[��H$�eqX4�������o�������������4��B�#��S�(}�w�z�M�vc4���������ku�yp��&���	\D�
Q`����Y&�ߕ³��n1jh�F � |k֬�v�Z���}���%�^*�tjrZ�d;;:l�<9L=lQ`��3�oF�2h� X��룵��QS:V���T0� o��m�"1�����a�8���
x�E!��а�Np �q�p,� �馛���t�b\��&�)������#�%��2(�C@Ri d�csK�L^�o�!���X��_'L�~}�EW� �Lr��j��I�+\�q?8�wu"�� ��''(<Ca�ڍ�x���y�D�����P%99z�z�A)�+e�rܐN�ǣgI~L�W�y8�Z�ƙ��1)óL9��C�.�.
,�aP{�r��c��=%H�!�E�(,M���Ć2����h��q���1�yE(?��˛2HA�����О/�nO�E�4�����k>��:d*�2�)2Me�aśW��F��`0��v-�������ql�c8�����X7:���y;�[YU���"@]��8�zLf�޼�*J���&J�RIڱ�cO�[�*���?�_��я�+G��$�͞�n��o��5M[.��N���"�
5Ey gp��ûhͺ����IIns�[�n�Tw�XBCC��˯��\x	{^Z�)R,K��N��ׯ_'._ �����<92"��뮻�6n�(�(J���˯�m�����N�/G��ˮԎTɼ9./�	h�o����_v��tw�*��T2tT|b�t���Fw�����<��ka��BW\q�������y�5}�J��&��-
x!{ ���P}#�X4�����lbժ~�̭���mq�!EjF��S^��
��O(���/U�&�k��b�2�z�r���x�����)�k�Jl�toMX͕
ܟy�z���B���I@���!j�xp�a�R�*�豟�3���84��=��p�.��w����_j��k��)B�Q�J2f��3�ju	��7@߃�n	=�Ri?O�|ܣmŎ{������HR�~��ՓwQa��g���0[��:���!F�c�R~�tC���p��FT�z`-�w�n�>���k[LB}�:Jj��<�m��B \V:l1�@6sn���,B� �]џd�� ���<��Q�+Je�E
@CV�JI�CU��ڏ٧1nP�d.��
.eךNQ{W���Ǌ�x$n�ʞ����dH=�t��^��[R\+Fx"�D�i�f���h�-��R�$K���2JǪ�N�FU^IMb��s���ɮ�{���X(�)@���7����{~�Njb@�΀�/�6���R�㶏����I#/�B�Z:(Mґ�#��7�K���OQ�9I<�����hrf��|͜_���x�%R4W.�Ӗ���@�zQ�`$%���HP��Ƣ:K�Q�_dX���0P%P�ntd���|�%�(���P�-��&��A;�ˋ�(O��Q�h�\��
�ׄ%��2x�e/t0,˼�f�ab�6�8�ny[X�Z�\�d���	�r��E(+a�"������q���9�d8��m��
�j�EP)G2�v��]���8��ԩO�����>X-莎N*rT���%��ˈp����� �̖H�b6M�<
����Ѷ��?O�s�0hoB!��{,���R1_����w}�֭]�����������'����_ �I�����R
�C�X�:۪�z�O�"/����K�{��/ЙpYuq��/N�.�}���tx.��e��C���p�e�'R���]����bO�4�3�C���>m&n�t��:�����jԯ
���=�X��b�p8��J��3N$[���(�k�r� ������C<��sj���T�t}�
v���b�k8z? �x��Ԇ)څ��kh
���#���|S�T��C�bq���5Q�� �h��e3YV��P������	���X�gݒoP�E�s]��іr��3蜘��$�T�����G���K��''��5U(H�f�m﹍f�W�ۉ�@[M:Aw���}?�j�lb�����f�R��V�T2jJ
Y�ϐ^�<?�,�I�h {�V��ޔ|G_��Z,��������:�*�P"�t�b�k�Z����?>�z#� �D���<	1��`����}�j�W��jRs�Z�:ihx��G�:��d�K��cr�Z{i/{q�Z��,R-�4^�Rs['���ttz���2Ś�{Q���LJ�R�r^�:[��o��oh���#'����z-��FO����d]W����[aa�-�WMBݰ(�[&6"���?3JE��Dd��5���������;BwXJ�&���s�G���9�������2�\5�h#~�� ��8���� Rd��6(��ª�Z�2�H��. ��2`���@L�����x�I�*7dy{�Ef؀S��U���vb�뷴������a୕&3�)"!+,&	����L���]�L���J������$���K�H���{t�7�w�v3�?)�Pmm���fn����J֭�о�������e���{�CW��J&Z��I��3��4oSMFHe,}u�|-�OZ�î��������V��e@���#��q��kĭN�T�QDPYdGSe�.��.)�Aw���b�7��g
xE��S�PL��/��mS�r<ى�y��>H"3����kGh�Ïs��h���xk+�3�&���I'(����X�9����J%Ds��u��С�d��ꖋ%��ׂ���`�+4�9���T��ɳ�CO4�*���u�������]����q`*T7�z�zv���=NO���x3E�6✊P�V/��,�/R�e� dO�}�vu�6�k/��˛,��fx}K��U3�*ʹLey�W�I�9�H�Q<��\��5�ß[�)xco}F�tq�>>twt���,���7�[O���m޶��n�B{��Qrn�P,�D�.��*���ҫ����)��O���Fk7o�D;um^G/+x�d����@�)����dy�b"��8��)����U���C����V�����}_��� t$�թ5����Q�R�o�e�W���x����T��)��TUDV�)��;e9�hI�u�I_�L1>�����Gw���0���hmZL����۷�y;��Df��c�4�zIɧ)�pd9_=p���^:�&��\�f̈
�{rr�4�]�Bc��`״��m��A5ӫ�&$��ק��XEu�V�9�ȣ�������i����pc����#`�e�(�O�2do��^#�Ë�m�4�30�%Ϗ�9dw|���Ȁ�R�!�QgC� .��W�X�F�I�
%{�ܲ����#�YO��!ҖeEOd������O\�*5At.�V� Z���SS��f���lNɃ��^rE�$ ��P�3v���ɺ!�z[����{��j,�}�>�̮m���	n���Y|N�b��~��'����?������U�i��	jkk����y�P��і�/�|>K/��}�p�4�R����O���y叏S_G3��%�+���pN+�$�\����Qˉ08P�=�hL���T	wZ���x;��a�� 	�?]���>_o$"E�Z���FE�v�l�~U�X&z���)��%ZH)�F�R�b�y׫���\c3Y���^!��󸩾y���r[�J�C�ٱ�f�'�6߇��9�39j��458F/>�M9Nk��i.7GV2F���ݶ�6]����9*�q������}�����vX��s����}�SoG=|�f�&�%���B�n�(��d�u��/\[8�U�G���&YPׯ����.���	�*p�U+$X��pO�Ŋ���ѓ�455�_y�����1��i4��V��+\���ʄ��?~>��
��⅓r5Io@�F�y�ћqN��]�&�5�w�p �>��@S��r�ڃ��F����h��*O)'��H��ó����d�t�o<ؔ��<YKK�������b�Ly��+2c�/X>\���"��.�[4���������ߥ��������)9�9ɸL�����-W\B����ԑA��L粴��h���h��U�����(�<|��`������Og�qN��%�s2�0�ߋ>����]��R��W��<�b���k�.����ʿ�^,�f�������/�ё&��}�U^2��ߔ��S(R{4���8��蓔��H���<QJ�4����5kh�Q�����&*{E*BV/`@<�cL����T�D�a�'Wp &+�
����b��	���\O'<��f@�}g��>�]�B���� ŇIVL�Y�dׯ[�T�˫�RL�k&�J����ԣm��_�[���F4���ۈs:d��hUb`~��`�"ً� C���0���B���  ���Q@�
l]T�I�W>� @/h�F@��X;��_�2�ZZZ���?���N����.ҐA3�P![�9ɶuƀW�#U� ��d��ZZe�9��+_�g��o�+����&'D5�\�)��BC�i�^�G7�q;��կSv|\lxWuv���l!+���(����-0�v}Q��BK����oW9�P�0<Lŗ�?hW$c�ȧ j���*{��t۬����H��ٚ�p�r���=�
-WN�~8�����5��s{2	��
Q�cE�_�FO��=/�ે�#���4�2ЭD"���L�]w5Y<!* +�N�4_'��E��W�Ux�x�a�e���Om�M||eQ$�*M��)�� Ǹ�g+d�m��$q�U-Nԕ��j��WԐ�ϣ?"�] Z8^u��O555ͨ��rޖ(nH�9�p�џ��v�ȏ-�Z8C'kD#�,� ��P4�U� �ZI-�\� O��m遽6�k�\N5�Ȳ2�9]ءvy��ʵ}[
?T�W���*7��#�7m��� �����x�	��m}��b��R���yv$s��3����SW�����&gg�W~�����i�;�駞f��JQ%H�L%�����t����*�%�b��m4��k��׿Co����L��P���0��n�"�^��`+����2���T*�)	��X#"�꒽i����)&�����*���:�넦$���R�d�ꊒN7GWv�
����|��n<x�1����V'f����������_b�ʟ����g�|�M���IS�<U��F2F9�b�PkG�ȿ�\��{�G}=������.����64\�r�"�i$�4���hY[zR<_m�C���K�{���
�-�ø�!r�y�_z�e��?���b�(�e[Y�}�DBQ�Z�p�-��V�i����Pbh�9�{�J����M�m[rl+=3�9����f��*�0fiO�����f*[a�k6���^`�,O@q1�?��� ���C��d1,B<��h�e@�V�~Yq��|Ƕ�K��@�A'6!|�o�������3��p&��)��:(@@�G�Je-
��0â2���|F���8�D�T��)Q�Fm�`N�g�Pă2���c�"u�k[�I�'n����أ�u�V:z�es�����D�u�z?�!z�+ߤ�����ŀ
'��������}=4Q*P�*S,��[Ff�RT��M������~~{ �U��]������O��5K��l�Yj��j��}�}�[��7rQ^P���zaj?u[�d��V���~��	����o ��*��|�H��Kh-!�&NR~ɲ�J^Mڂ� ����hs%B�<�8������K�a�����Ic�<����Q�ﱡ�y1����	��ESi�df)��D9��?�O%���q1Հ]��*kY��k�`B[љ����[�C]W+\W�w�$4�Z�Ke��Q����Vk"橍�3���+�J7�V¢���3�C4�A@y�1>3>1N7n�{����~&�������m�m����D4"nv���E �@O�K����5�_��7�hסWg94���˶�2��LC֬oP4 �9g�t�l�(D�;�-��R=��Am�����B[C<��t�Y�7�T-6���IZ}OW/�J��f)� o�q�h�:�ev��h��5Uy@;����rrrb'6�({cZ�QHe��bY#Ho��v�z���4��rͨ�̐��T{kM����~�g���<?1D=}�493+�*��D�fgiͅ��=<���_���)���|&'��}_���{�-������H�{�ixd�b���)x��˕�5*p�Wf)������^��WyfW���}�g~�f5@��(O>#|_Derx��Ľ�Rqt�z�Md�<�x��;�OC�]w��Tb@�*��ꔟ�c���6�4�idb��[[�`�k_���v�ȴ��1�.<���,��&�gC��84:f2�5�^�� P�ad��y�(��>�s�E��3%�=m+�:>_�Z��u4uK�&4�ey��Z�}�s��͊����h��ۈs:LfWt$1@��Ț%��d�2E�1�Q
�zڕ���|���yv(KrxIq�+<W|--�XU�Z[q�� 4�u� ,fC$��Rk[�g[ZZ�05=mc���h���R`Q�������KU�Qa��d�ؐ�%���x$J_�ڿ�g?}�¯~���t��[Z%C'���iJ'�4��|z��У����O�\Yfz�ʳ3�ݯ|����wҪ�^���f��RP�d_�?O���/ܔn����e��T
Ѫԙ���`��&#&-� �,(�"�VʊP����'��ӻ�����ߗ���$��|��je�Cb�������2��܇���2y��W�F#C�Ԝ�����Hu9���b�0�,dnaJR�*B�z���=�+`�jlr���W_�����.8��}�$��y��+kvG��qsT�*\�m�Z ��ݲ�h��� ��8���"3R�jU� ����898���a��DȂ5+2�<�X�⬩A�s�*�rU�3�ܕ*^���ɨb0mֺ%g,U���}���s��n�1� �Š�p�˒R��diz�rQ����Hsp���ʊ)'6_2��R��n�H��ψ��G������AL([�R���Ƨg�\)Ўk���|��ߢ��YZ��K��C4���o��e���w��Mh&�����uŒ=_'������ ��t*�ؕ>c ����5l����R�_76��f��n��(�|�$�N�/�B��C��۩��S�/R�)E�]��w���L�T��^��X�N�L�q)Ο��r)W���Nz��鱇��k��Љcܞ*�<aj�ёJD[�G9 Eg ��&�~`��Գϋ|>�m�]�"����ݼe�Ȇ���7X�爫�Q��x��V����������ݠ4��(���`���U�\O(&m)P~�T|WY�s�P��j;���UKϞ_�쭧�я�w��T��V���V|F�ɋA�F��SW�GD�-%n�+EsQ��7(��pL;�{?���Zȼ�§�d	�$a5�N\H�+e?�g��B���X�h������z0>�(��d�f�-�YV;"
}�O��҉4���?A��#xm*����ԜN���]E��G��{t��	jmi��h�$?z�tE�H}��PGW�=qH�Nv4��[�R������Dܘ�:-�J�ڷK���V6`�>lS���DLMl5�r���BF�2Ŗ:�Zw9 �(,�ֱvH�H&����`k=�C
/�d���ExR�bE��#/{�N=A��Y�d'���lm��U��C�)��C�ǥR��g����2�v������'���w}���І�Ut��!��;���\!OY�+-�U���	��:&K��ԫSHs��+m�昴rL�j�mY�}�]1S�D޳d�U!��V�Z��<L�t����?�������̌Ȕ�.�{nr
��P������>n�r겺u��泍hě-���| sa�������@S���s���� k�2cV�����2�Ė��Z�CVTۇ$�]���OdW�Υp��������ook��hS���L&b�2kkj���Ų���T�Cj�"����ܵ��|.O]�4����K��O��O(� �m7�(���3~,��6����&�i��;��}�v�hg�f�����O�w����'�'K��ۻi���+d��:�l�/H��#�1�EbUG+}>u����:?��p%ӚƁ�(��B�]����"ۯ�*m������=�/-N��=��y��|�ē��1zm�:��eʌNR+O>bPG��޺���n|�M���s���w�'9Y�o��1��~�yze���� 7;3M��)��4��F��m�x")xg#�%V�g3`R�*�p��<�Я��cLJ������z׻�	�8S��8�2�`Rb �Ei�����h�J� ��8��pӌ"� NZ\�I��7X/���Ǫ�Zb�m���D��MI-�b8A�{���W,��x����z[���y"A�}}{'&'���oƀ�+�n�d�kϣ��`�p�2���z9*UCg���u6���S�y��e(O2�ɋI@�W��~�W�K_���y!�D�| ��etv�ڢI��+��������(` ?[i�������_B\%�'��Ԕ��l���rfs�׍�3T6(tB�o��f��ʂiqO��(��.l _y!�P�]G�6}���	�e��gSp�ٿS� c99��mI�O�'��e�Pb����>���o�P���4����4��wJA���	j�2@S��n��T`�E��d���Q�{+� ��ϋ{����>G�L�n����
�Y����'�<0��k����؂e�/�`�t�C}gE���-�|¤�Zݤ
c��/�P��٩iZ�v]���~�';;;''�&xb���28́L�]�����_M|��|�k5����1��m�)��i����w�L���X�f6�TA�f�4�H��`�犒��R7�d,��1�[𭏈a���Bכon*A`��v�y�٣���kkk+tvt��D"�ߋŢ�ϕJyJE�*3z�ﳝ᭗iB��k�L�gw�'NNN⛒�C��Z]�m�k��K�k�.jij�H9B�\��(���J��d2�w�f��/|���^z�0���R~.+��O<GO?�m}�E�q�6j�h����ޒζ�eq\q�q�V�u3���T�����H��Vذ�}]�:	gX�t�MJ&ͫi��^�U�f�u��8c𠏸:	Y����7*���*dx���;���b�����Үv|�ċ��}����X��::�P�\\@���\S�����d��i.�S�w�^a�M%����ϊaI>����E�^|I	r����QZ7�`wnZ�R
�oHfg�du&���t'�K��%�L8�nZ�f�ڷ)j����k�n~�����ɉq�b 㿣�1��
	���jS(vg)%q�᳡1���Ù�X({�Ԇ�g�{���}n�3/jZ� N	�.�=Aؒ�#�W����������8��rXu�	���B./U��DR,9�����B�T*�~'���8���V$k���-���ps��v����d8(�DWS�z�L"��h����}5��Q"��TYW2xF�*�h�y�O�!C�"˞���RYYu�t��Y
��8�X<�q�|?�˧�m+ɀ$�Ɋ{�>�h�/��6���）����nz�t�� _��p4�h@����e(ho��~�?���v7��Y�2 mѧ��qzef���^r�����M�T^��CN,B�rY���h�_	�9�����˨Za&N_q�=)��M!�\ QOe�M+9x�Z_4P�A%]��~�&kN���J��W���S*!8�hT�����{a�.0W�9����G>���o_U��J)	X��y��O��O
=S�/�]/P��u1؍��+<a�t��d�bM����Fv:��r)�`���ϕ���-����c�o뤱�1z橧i���b,�73K�8�e�a�!��U�������ߡԀ��f���岢d��W��J��p��Xh�����gn��O;u����~[�*�Y��H��V\�W�����=><H�k�~�w~��gʥ��g��D��T�d�Qo�¾OQ?��*Y�Z۩�-��^���R?��VT�Y��V���=�Os�9��F4��F�C���ּ��&���z�o� �� @IZ`�r�26ЅE��x��;[D�S[j��������'�-uB��X��<ZS���e�����l�gx�V̍�&_;�)����=��y-��D{yb G���n����cǎ
 �J��� �@ٜ��]����_��_����ߦ�������I
��9
b0��6�A��)��?�ں~==r�w����ԑh�}{t�=412J׿�X?@9��9��)�b ,����^�A�Mq�6�`Kk�ҭ�&��e�Aep�+����v@���jA�ڄ*��C�T5��i}���HP���B��/������A�9��%u�mQ��Թ�e���؁���.�t�hQ�/�˯�"�N��������Ѫ�K}-�D�(M�5���u��k�o�z"u��2,9w�'K��K���20�li���a���^:��A�X�˸�IfRm�yʤ<{d�yB�L���e��ɘ�iH�N�y���o���g@�}�MDTџ���Dn�*��+"��B�]{6���W�|����>���g-�i��j��^�NV���4a/��)���{g�a��6~�ƿF��h �F��a���:S)� �+����j�-�=T�۪!��P�4�]��ә�4C}�}�8XQ�g�<]4�,q �M �ֶ6�ƍ��������	�N2rV���7'2�S��=��?����r��]{��hӦ�4=7+6d��a��\)t��u����Ƨ������^���~�"���>��t���� Ȋ��Λ����.������T+SY��f(���:��'v��b�z��i-d)Ʃ���'f#Ġ�+Wȓ����MX�Ws*UUo�t��Y�7��	l)�*�V��F��8�b�Ae��'1*�ߖ�:P� C����^X� ���S	���U]I�52)0�Z`��ѵ��hL&Ȩ"S����� x�IP9W�R�GSG�О}4yl�6��(;7G٨-F	���^���֮��۷R����ʼmP�0����"��PoW7����/�f���(4 ��2Y�f���1��/\q@V�������*t���Nh�	�_�ւ]s_�I}���Ả��67`W�M�j�/���������]6��|����LF�=��(08�J�g�Sk��H�6�KE�6����,/�a�g~�l�Ԫ��η��D/��u�<� Z�KW;���S݆�eO�d��^S�m�ĪZ���?~���驫@�P* �st���n�����.�v��T��{dd�o^ /s��֯�f��f�]�ٜ�P@�����4<:L��o?G	^#�C��@:?5Kc��-xy?uo\M���?�o�_��G���v�a ������}��g_�K���:V�Ք��_��r�2�
9� ��fL _Q��;WG��p* �@v�sW�^��|۶�Enu�WQ<wVT���I�ڇ/T�����0������kn�U髞�3Z!#�|]!P�Z��/4-}�w����� ���R<�hpik3	�|�L���pO�C�>H��Q��D_��
قh(ϔKb�ۿ~�6]��bm�T�Gi���HS��\��R0�"O"&U�l����K��J���(a9����B�RN��q7e�(l����_�i�<��T*M��m"��Ie����@o-�=^W<��j����`W>��wM�$Y����q����?�����C�'y����+%]g�6��){9�w#�c�ۈj,��(�A�u��Z
[¥�>䅗� �,#:CkJ�R-����t#� �,3�����b����4&˭0� �V��Y�tm-}�P������ʔ7n���|_?t�� �_�	�
�H4�(�8�v�/���W�ݭץ]��x��Ā���.`������d�:;:�Vw��~�(�'zɼ�$�R2N�� ���0}�3���[Σ�Cck���i��R��>�s��H�M?��y�Nz�{Q��!�K����T"Is�c��/�E�/�T��7l�J�m�487������ɉEQ'Jy>V �ńż Eh+mǪ)�v��_�? ��k�U�t�k��UzϵקV!��!`K�yz�����qH�ѥ�)�4M�~�ͶԲ��h�@��(���9��r�H�|��W�o�=�,����Hnx�^~�%:��A��eh����)��!N�X�Z׭��uvw�Oіe�Q��fTSy�o��=���A���������}��������eP@��n��Fx���W?������� I��Y���r)4����WK�9����=�+��Ү����.^p�+k�F�g0!��T���z��'�+�{�[���|�y)�f�U���sR¾�l��3+�kD#��� ��8�B�*�Ю��`��}ZlIRV&#��$�Va�H�	�7P�Y�����a��ޕ�DPN]յ�ge���q{��#������U�N�������A�u�Y��� ��d��I��g�;91I�C�t��qhө��.�&vt@HF���>:t�0=�����8}��oZ�������k)��QɫPsw'��v�����E�\L�ǽ�ă���y�2���-t^z�)�81L3ãԿm#�� �)Aӕ_S�Ɇ���k�>"��D� Kq$=�^6J!�[@��R�5O-�[�a-c����`�t�2�P�~Ty�@�b���I�m�t T�d�d+*��q�t�2<]U��d���)	7Ai'F��in�!;6H���g�[�J6/F9���=�d[����G]��S������g�}q ����d]{:�(������3�<C���_�0Q�/���j�8Y!�<cӫ� O�%�@[�����-n�e�y_�H�^,z50Zd��G���I�<�3؜G���{+��$�o�v�O|��K�Rc�ܖ�*��ۍn#���xq΅��R5 ��,@���t�z�&c��è�aEњ���(
����� նt1[DF"Q�2ȵ���[�TB�˸�s���Ń�gy����.!���X�]#+4/�j-X�/��βjB�Omm���.�ޗ^z������8_p4&&&B���bt�$5��H�nt��mo/��������>��OӅ\�ۚd U����_�T{y2A��Z{�����;��ޯ�CG����AZ�z�-T�����Ӊcǩe�_�z֭��>��dY���ƣ�pnKX��������ca\�F�K@�B��P�e!{�%��-ͩ�'dS}�Q�d�����.��l�_,��_��#��(�|�[&`�"����hsu!�;71NQ�Rv��-����4x�U:������T*z�$Ҕh�6����q�����/����	bq��e���2 �dѹ5%C�����۷��z�):r�JI��m/�U���W3�ՈJ.�p�M�w�>��i���� 4� ��Vh�����0nj��
H(��?���	���4}�'>0z�Uo���Bٗ�#H�X��Р,4��?���s����k�����T$��W !%�����8����R�8�6�[��%ٮj�W��,C[��yQop���xw����e�|O@9@��Uu'��������������l�/�BeyΌ�[��z��>~��2P}���J�����pq.���"CUu �ڧJh�sKK��!�(<��Cs��ӳT���ﾝ�uۭ����m۾�F'�¿E�0�/RKO��SEr�Q� F=�bI����3�r(Ə��B&O�� ����/���o�B--ZrE��*";�R���+iU�*Z���V���}���+�_[�Z53�k�9����_��W�0�;�}��$.Zv�x�v�1���{�S�P�T�jR\^��D�����G^�@���������Qj�&hms'��g�7�����������;�S�yk)��Fen�i�s�9�ٵ)
7��RY�y'N�Ҟ�{���7�n6�$�܈���l�V�� ��P(ݦ��@a�砀��J��\�@�x�F[Ds��c%J��s��}�̮�?���|�(�l�������O���d2�1'���u�*��/c-`�c5�ш��xϡ0�o�$��g�=�个t�SU��'�F�hɒ-c�8Ȥ���Yc��{D�s�o�KX����޲���,`�ŀYL0���g��aFa�&O�T�?߹u��kBK��]ǿ�h��+ܺ����~����Զ��{��^ʨ�M���Z�TTj]� m��%��T��?G����i�5���,�d��v5He���8R�9%��u� d�yN���J�i��*q$�l��^�	�����#r%�hx��.�B�P�vxx8�*l�a3L���J�]Q}�]�EKU|�I���[�6ލfF_K�u�(��d�|> 
h�d2A�z/�������ln�KTm�	h��
�
0�#k' �\��]��� >�.^��U[,&<е����n�)=�ȃ���|�^�W0��DSI��G�9��HP5�Ha[d��|�%��Ï���Dy�jS|�� ��*��!ع��>�\j��xG+��NQGO'uD��Ie@%b(�t���$(h`� �|�0>�X�� �j�L��F�"S��?Ȋ�o	*��Q
����`B��6��c\�0�ɚ�8Ⱦʢ�Z��เ˜e["�;���b���7BT��H�p��z�v=����O���m��m(a)^;��*v�Ƌ�]��κ��Աr1M�e*%�4��PنDR��r.+ϋXg���ve���{�:����4&�4	]l/텯?�r�U�P�ު㵲v�!�ߕ*T�~����|^d����|^��	o��7H?�}���+n�'��x��]!�<��:��VCІ���I�(i�CGӫ^��a�@����=>5��YD��L:��W�w2��
)%�zȿ��s�zMW+�D⏛"���=�⩾b5�N���d& j�\S6���.��pM��ltx�����P(l�]v<��r<��LeC�}TB�̿�dɒ�MLNndm%�T=)rH�Vh�,�n��2�-�!��T�>|xV�Rx�$+�z�j+�)�= _�
٫�����7��~y�m��k�H�]�؀����<�5�b��T��Qe2Nk.8�VmXO�Gh�ȰpEͪR6p�e������/Z���zW.��kVR<����h,,����0 �h��F�
NU�͊b�P��T%I'K���� �q�^J��7��3R2t�B��k �L�l��������me��
i��E�֘�+����qM�|T
H�z��p;��F�68@;�&E~�t�Z��OQ�An��FD��[�t�JZ��J֮�����nIP!7�@�H�dL�����E�hmK�Vwg7�q����`P��C��%m"�f!Ugp�wB�X�W�E�\K��� �mc��l)90�l���.8� ����ֶ�c2�Q���Ź=�e=::F�H�����쟻��G�L���0�	L� (|.>�!�{MO� ��#D x�xZ�����oU�W+�p�[0B�r��D��������W~薅W�rN������f�;�nݺ�f���SSS��2��,[��|f���z�p��3ɳ	�#;���.��Fcy�o�l���ɚ��c7T���. �mi
�$pI�A]{k����h���o������?Ц�73�5)��j�J����E��hrt�������nY����;vS�t�P$�{|���>4D�x��:iѲ%Թx!�e��a%��c	����N��|�9��f�5�HT�	cSM��w*�4��E�Y^XT��	)PdUUzP8��a���'����E�����G��EeaAؠ�T;Y���>��kA��
����6�Ѯ��������Sex�bԣI������P��a���gQ{o��[�Q*0.r����!����qZ���֏�Q���7w��n��b���s*�U2u�U�x�x) ��梟��j	�����O6�rhzk�d7��h�b��5$��Y�QY[��3iz�5o޼y�u|�v&�U�ז�5�J�i���w��ނ�� ��
M/P&�2��dyI�`Q���3< O �QS��Nn�gyEG�q�z����+og y��ؘ��`w���#$dt��Z�	@���U�V��Ď;�M����?~#jK�罒pZ�XO$iU��8�' /����$�[�R�}ÌQv=���ʫ���W�ʷ���f�``�E���C�����ZE�C#�q�Զnm=m����y�ؽ_��Q��������s��=460L�w���NZ���b-)�a ��l�֖8���M�*!�
&lrM%f���3��@�.V�c2G��(E�A��!@N
��咢�hN0\�@��lC�|�V	�)3"��p+�MNSi:G�r��w�v:���
%̨P�=.�Ӵ�w�����e��Z t�8�V�����m���4U��#FDL<Z�)�g�c���{�\{zz�z���� �x�馛n���1�4tQg{;���;Q���}OVh�@dye����^����Y����	^�>V�׬k��M�X��Mt�'Ae����V��/��K��Xɥ%S)*����xإ��7� �H�7�'5�	���U�'���q�^�����V���V�ՠ�����Ga��H��kN��RT;�&�=F�l@g�\v:�T&�ܔd�Y8���942|�v-I�)K>c׎9�匙��f�3#�PP�+Y�$�lE�ha��|�r���P�݆㹧Y�d �[�>mY�uQ��@����$Hg� �Ov��S��^�pD��-�}�S��������7�s�s��_O۰�
�"��NP���R=�4��wz:Cm=mt��Rab��?��v<�(�Ǩ�@�\�0�Q�3�L���;�R4�`໘,���=d%�<Z��L�h���d2J=�-r~S�i 0A�?�����jY>� G�L���]p�n�T���f���	ro��˙6�ZCJ��O�'��4M���q�ML����T��F08�Q�6��-Rٲ)� ?�h��ӈJ�DH�.\��6����W.�hg2T4*T(ɊE��P))1��׭^#J1~Ag;��?�����44<�`�ȓ�.)J+�f��_��a7d���4�wG�a�
C����"�E��7y����4�����T�5i3oT}�ܚE�O���gg6�6��Xs(��
��� a��YKg��l��W\uh�ik�ɓ�X.�5,e-*j2S�f�,m����:ݲ�DA�̍ ���P�]�Ru܁���Y_f�`e�5v�C��u確��LF2��m{�b�����.�a�MX�vvt�Z�f��C��K&2�b~ �f��דJƬZ�'^�x1M0�ΤӒ��9��� ��0?�֮VU�(A+l������A�F�lN�u�Ci���x�"��g���u]y�+�-oy�X��A �:�;[)W)����o+�P� �F�V\|��r&����G���}�����b�$�T �����Q�<:J��=n�-Em]��.��j�����$S̠��q;�������E?i�έ "G~B�8e�ކ	�~������$;�H�0��
8_`�;Ϳ������8��R:K�LN$�/�!L#�t�|��G���� �+Իz�~�Y��jOQ��ReP��|�G�� �>1)����V1��y2���A���^��o�={�奵5E�v<!(�BgIF�R����Ҟ>��9�8¿��U�yB�VJb��}W��*��'���(�ԙe mL@�w��[����k^��f��	� ϰc3�jq)��z���<��EA�| � �ҡh�����L��)7ˋA=2T���WU�����*���4�a6p����2pq�ע��f�kI(�w"� ���Z��s�vﹺ���� �X���68�4k6��Β�J�]�����|�ή.}{��72m��sI$�T`�e�\_F��ڦ�3 X�Wv�f-륏��5�C1����p�dP��
�-q�dS����o��qӭ��7\Co}�;i��N�NMN��m8�MOQ>T03RK��sV.�s��iz�w����C���B1���� �ltfd�&G��5�'�B}Yo�0��-���8��J���,,O��x*&�(�L~�"%�z!�Vm�@Dn�7\�cO��M
�>r�0���}}�;�&t�`�uhI'�1�B{E�9��)�Z[;-�s)1:�.�c�"Z���v�w6��&)�Q�Z%
����qJ�
���������.�:͠{bl���ߠ�n��b�?���P�(iz�(}�%����d��ɦ�p��=gE�����/�qW3�d
`����2�;)��3x�ȶ��׊P�ꮌPd���>��_�P"�q�R��1��ERL����*IE��:�#"�y# �A�R�J���t��Y^���:�,��C] ��t��.8�%#l9�z���ȱ����(7+7{�x�O��l}�Ro�m�U��3CV�5�*����+V��n߾}��� Xr�8͔��lר�8��L��XB]�t)��'�� 7W18da �aU�>�I��]%�����978ё�e���ͥRT$�:26*��q�a3D!�@�#��/|�n��fz�k�'���o�ŋ:hhl��siu>!�t�&(��2<:JZ���7�}��_H��Hv���M��F��*d��+�Kk�e�D4N� ?]�"_'8��|��"����ۋ�9| �����;���)`��hI�0`� D���c�(0����wU�p�����v.��T�,LϹ��C���\�C��,��Z�e�Z}��Խ���X�F��:STǵ�4pU�[��=�+�~��l�j�c��_�v3��Gߥh�d�Z/��s�� ��"Q�ذ�n�����`�u����&�w��ն*ӛjk%X�"��$)W��T~[�]M�˶�߯�	��6�(R����5�3/��Ͷ��s<'q� �.�I$��z�θ\�Z����r�U~<��� C��=�{
�SA��x�љ_�y�X}Fj5��ڧ}.�I�P�=�5�m�Y����v��)bրEU@*�p�	c
�*�\Z�S2��P!A�v��VX�Ԛ��#��ɲď�'p�p�u����c�>�֣G�.�̏�7@�*� �nG�.u��s�52�6��9Si��xB@�,��g tV�^)�>x� ;�N?�&�,���R�u��2��JW�l+�
]��	���^����BZ"�}˽(�B����2ɩ�T�X&U>#��x%�������]������'��-Ϧ5+W��T����e �H�"�V�.�)��'��`�"b�pƊŴl��>:B#C4x�=tD����2���̕
9���!J�"��GQu�{����7�V�
�"��ݥ8I<� �P���ɀŎh_���t�RVBګ�'l:܇��^(�R�k%b�����b����B��k�.��p{�����B��EwN4E���WD6F6�O(0��> �m�m455;l�o۶�~����;~M�Q���jW�j��(�lV�����5��<�u@�B�&����ŭ�%&Z�wF�ud4�������	˿
|��1&_ ��>��Kc( X�Q��L�,w�H��/�.<�K�����cD��p�_羃�S�'c�N)���k��������NGQ����ŵ�wk���)Q��q�%+3���/"S�N���N��ԇ���p4�Yl:�`yO<��S;�ƯXMC�Vgfc�$ë�ܬ �qj*��AE�F�%iw(�p7<T
�nk�7��h�VӶQU��ZX����?�K���/��h�B�_�Պ��d5�����D`W�R�= <��Y�n�(z�%�CNT�\�>W�<���UePZ��i�yRR6�z�O5�R�-���*XD������]�2����ut���ix�(����^9:E��V�=d�Qv����A_��Թd-ް��(��Vibx�������622Y*�roQ0W`�L�k�F�ֵ
r��jYLSLe�2�IF%��T:L�\�+�(3X�*Ud�0!``m�O��A���)��F�T��l�Lm�]�.a��;Z��7FUF9�({+��)�ٜ�X<AE+#Z��J-�8������?��ﺛ�8&o�`Ae&��u�$�a��B��%K
�`V���IU�J_�t��PJ ]�}կQZ
�h�l��sfH��k�:2��kT��|!+�h�~񜅢J�������?�g}&�/� ���Y�������^[����q��� .�L� ��
U��z�J��(�B��!]q-!�����d��!�?_�V\�k�z�u�㷫��VU�����F���� ��g�}�7�����{w��`�2@���l�(���N���X8�b�ZQ ���E$�P��C3Р]��@3�.�X�&Cf֋=�V��Ư���)�}�ܔ]�ɱ#�ӗ��e�ֿ^O/z����׾��<kau�ŀd"Dmq}��	1�p�S<���p�K�i��.Z��3(��^�0��G�Pfj����	ב�r�
ʆ(>6x�4d,�><�½%�ͦ,�n#9�6��2��|)�@ˤ��jik�	Y��P8�%+�S[G;u�.��dE#���T�Wx�T
Ǩ����Z�rIؒj�ud�jm�B!O��I���Գ���R-�O�_��6������ `\�m�7���� Pӓ��=��Ď�������������YXP�`�P�g��"�O�;C��2�DX�0�wJ��.�����?��Q<�>>	���.��=���j�?����}?`�?� �U l穰D�V�7��]xA�_QAgqC7ej�>`,���L�3LU����B
D�z���/�s�UQ^8�!C	^!2Gn���K.�Ԯ�;��\*����fy�~ߣ�U4��/Yց��kǠ�5 ā�#Ri�e��>+�b��γ;�#��3� ��K+����������
s��F�dY�?��XX/�����&���N[�����o��������
�ӦMgP�A�`bl��0@�ENYP�"I�zF�<��d�Bf֡��~'Z:��%.��w�� ^�Q�yd�
�9t0����W_�Mh�78��BI��&c���P
 o�d�2��*s?�EqFDe{A���a��+T�"�1p�K|/�%����d����v-��w1�1��;�F��z�G��J���3�4�*�
r�:��)�N7���"O�	��҂�+����� ^?��/�����q���y%��&������U�d")4!��

`�`�w���A�=��|:15m���c���7�<	>%�H�٘!ѱe��"�z�7�'5f~)��%��a����W���[(bפ�j�70x�����w-���Z1�.�ҠL�7�2Ĥ��
$�b3��[�/�aq�Կ\�!C�u
�
E����:k�{���-�d�����-U%�d�y�]kQd�n�9�ׂ��]��֬YC}}}Be���-z���k� �o�]U�׷G�̿������~�a_�}�u��j��q%ܖ|^nQ�i�L�ѣ�Ԓj���)��S<�����}#���O\t!��ˮ�+����o?��2*��m���~r�9ܣZo�bS��5ڑ�r��~b�dT�5!z�(>+1(jk[G��ꚋE�6����Wo���	�+�K�v���u������i���u��
�Ȭl�3��J��ɶyaQ$�x�|�Q�:r�:;���{��!z��?�o~�z���)���s'��<��QY=�糲�ђT�h#[�҆���t�Rt��@��f�eO3C{�����E����L��⚹�>��F�*��E��P�5 ���i
�^��z�9G����	D5$td��]�6��׵
VIE��}E��Z����,@���/��W+C�wu�9�:Hk֮u�yӛ>�Ng�pi,�
"�V*cR�9�j�2ս�Ɍ����8|���U&q�)޴d�=�?AD x�x�DMj?�- �Z5]'�iy���%y�6Pk�A�vj�^�ؠ���¼��S�Pfp�����``-g����;�����~�w�ޔP(��]�}�1d?�e}�nOO��+,�b�G�<4x��t
�q�ug�&>!�n.��h۝��m� H3ɹ����֡2�0�K�dA-����ｇ�����O}���E��կ~m9�|2��d[A�V4�l���%�	��⌞L���2���*����8a����E[Z���ӵIS�mC�q����#(�\�(^s��-�oŹp���� hQ8��)�l'�3@ �T�n*�
��ɦ)�H�Մ	o��;~M���wt���2>��
�Z�D���s�����	9'LyMK�s��5F0��7�N�pc9�bϫ�����*N�.:�ۆq'��9ÿa��;�U�:Q.�j`W��lN1p���#��ja���#�I�U(�q��?�{���^Y�d�#ӹ�@r�q�rI�6=�AB1�E�d�퓣*D�� oO����*�㨭�V�W;&��o2�o}u�%FST! |�fn=�Z��u�,|���Z=�� 8>1�tuw�à�����Wf2Y�Pȹ��!˰d�l&,�t���r��q�pp��mO����Б��D�0o~P��v5�}2Cg���/{���>����@N�!S��X����J&���W��9���(_�u+]��ѕW^E�d��zZ�����Ng3����ۢ�6D��x(��0������],&�R�&@*|L'�4~�!��H�S����
y"Va�����C�J @���a�"j���Q#��9�����Gk"����A�޽�衇�;n���q*e����C2U`*��*�J��)~="���@�hS ��.�VlC���'IVkWK׷:�����d�����\ev-�>�J _/�M��dQx	��dy�c��E6[��\B�v��fX�̊�⌕���ʑd[Mi�'���~������N[{+M���jI�ѱq�z��Γ'��B#ܲ�2mAıG x�xڇ���[��39�����"�Z_�V�lR&j`5����K�We�uD~ht|\��<��7l�x_��o��Sap�L&�R�J1��Q#��8����C�_��1 υ�{xhXܜ:����R���9�Ɨ���U�����d�׵N��TR��d)�©-X=�Vi��(�G~������^2��z�9�~�Fں�b�]��V�Z��(/� �l�R*�F-IJ�%)��R!��0�ݮ�nY$1ȩ �B5�LLb@�eP^��B&�a�U�R"��$�P�e��X(<�E8���|�qNy�����}�N�_���;(���0ZGΛ���)���e�N�F 74b3�iE��g�����+��,��Ҥ��$�2]�k��_�`w�ϓb؊P����g�>�sdfU�eU��{	I�%Kzi��^Z��4Z��Kglڤ�\��퐩�9ˮݻh�����N��f�-<��3?K�xB�h6�K��G?�P'��S]9>9����I���P�i��)�懻O�4� �� � �Ԙ���g[W�s���x��Qê� 2h�R}y�6h�FP�_)����T�}-*d;�9��Z�E8���БDD�I� ?�9z
WkV����5+ہ�(f<�㉨�)]<H�|�Y�q��\\2wCC��5�)����2p�"C��4�H�˨��&�W%�pi�z�:3��G����-��%e�1-��aQ��]p+��i*�0{��oFs�f��~y��g����vWC`��+����N$~D8Q_*�@����1~�%�������ٍ��f�F��Z� x����U��.�e˖���i��v���� ����%��2�p-J�xK��Bm���PYr���e���R6��r�&2׹t�F��Y���G{���o�ѣC�3"��Q�r^q}�pcaS�ť�A��yR�_q�.P��E&�?A@� oGn۩����j�����8�3�3ǻJ�Y��E��f�]�W����j�O�U�/�-�鯱DRVHb�A�ܢ�|>'�ikg �hm9�<��s�Cؕ��S�L��D�y�|@	�`?����;�St������R�D+���D<)��ѱ�2�:���?{�e�H��������	Y"���H����8�K���BCu�Uio�<
3�v��>��籉SǓ'�5'� �3��).��:d���ԥ�4�fDCV�����!2Dn�I/}�e׺#�Q�����r%8�x��8�ί��bQimm��ƍ?���vtt
(�؅�~*\G�S��7�9 #�/���'d����b��N�]u
�=�HQ#�!����b"��m{��������i�	��َ@n�>H7�*{�+��k�]�;W2j`�󺣖���E[�a$1<�h��O~�G��_�� ^�u/��N?�z-��˗QG{ߣNn����Fî�E21�Zu@�Ng  �B'@V�'fG������~衇Ā`C;yjD�'�Đ��E.|g��4�1��k�S����������FLs���t�Ec^��z{6n��Z���>�g��OC�XYppet/���6��/y]t��z���=��х�(�-����X��G~61X~��^G����w�A۷o]I�/�:t���o�u�r��誏|�#�������6LD�����"�����7�<�D � �֡ᑉԚ�"�e�3�r1���B�����[ə�j������}״�Ui��9"��\=�rw�K{�\�u�����#���ĸ�C C
���C5z&��bh�nX���oXOg�q�ط��)��L��q�� �� p՚lcP��;v�#�<*�B � \�7/R�7��l�k�+���&��5 ,3'G2����C�!q\�Z������wg"E�H�*�gx� ��lP<��RY�� �'����Aouu-��TJ&)xj �B+��E���!6����
 �	x��xq`�,���R�@&�qT��#���Z-�;`-�=�˙�
5�{�	���#�5�lﾎ!tfW+7�'�z�@�׎�:20 ����N���X��%`��[�KW_}5]p�����~G����c�*�l6V�ܷWW=����LNѪ����Σ���n��V��7�A�me4�T:-�_��WR�?�����������p�}��L9;�(� �8� oO�P[���W]�VK��V�س�l�xkK�V�6��5���c�Hͮq�_4YfTʻ�1�l�:>6� &,T�{R-��	����gn��=�yt�E�Y��RRJn���&��_dq�Y��8�f��ſ��<�w�}t��n��:(�]���c��j�{L�6���и���C��ym��oӀ�DT��^a0
�&p��R�etvR����]�=b�D�b��w��&�ģ�0ܷ�LW��^�z��+�"��`�7#_�%�(�e2�����cQ�� $�#Jʫ��j����5�t"���	��se�E'�!�����dx]#=1���MLL`�X�D�a�,!s�.�L&�hgU�f׬��\`b������ئ�"�
�0q��q�/^Loy�[��o~3}��_�o�ے}�3���Eã#�����3s���>�ɿ�lGkky�'�^�5�3)C���$#� �xb � �R������:zI��.E���n�*PA L��(�TA�h�͸! 8E�C���%3�D���i�	|>T42h�K��T|���_���e��XX�P���}��]Ʈ��D6J+9 ��3J�\D�^z)�_��V�\N]�]�e�5~�K���E,������J���֋��ƍ����뷴w�^�
Ɛ�G���3؊���r�Ԧs��"���x��\�c�������M�^�k<0�3���:X��S�e�r$M	�[T-+w8�*�lҷ���pD�����5TA`��\oUq&���u��Yhܫ8�4okI2�m�Qp�����^Gk��k|j���3�\h�R#(Հיl��,�3S�`6�+ ԇ�0��׳�;��`�w��\r�.ح�&�t{#jz*��H,/nf��mb㋉�g?�~^6�4�J� �62֪=m� z��f2c����C�]�ް�U��k�.1u�D|�����W����������	5Ž��o���{�뮟��K^�`G�ũT��%�k���`�fN��ķ��	D-��3* ,uf�F]p����*t��2A0]�Q%�� WV[��@��F���@Z���1ؔ�l��<���7NNLPraܹҢ�կ~�N;�4D��v�v���|�&��2�j�C�1�-��t`�7\�A{Ѣ���+(t�a�Ν�'�'(�͈)�'�	��|�_�w'����ڦVi�����m7�ZV�����)�"���,)\���Гd��F�J��f��^&m
��k)���5��nA�B���**җD�U��l��ǘ�ϴ�������H�p6�i�~�� !��"xf{������M�����'�����Rtd�� Zp����w
���VЂ�F�d�cbr���dM�ֻ�3[� 0� ݪ�q?�����!Y}���b�x�x��Y�袋����6���]�;����77�e�͐�k��?�� �x&E x�xF�,E�����PB1 ��$�B/Sq���mm_
������Ȫ(�k��8����2��A�ڵk���m�v����_��k�W���G�����R����aJ�`���%��XUڊ#�d���D2&?�����vw�/�M�h���b� >p������	MM �L`��sz�ʉ���yg3��/j���OR6��b<P)�cX.`5��h:J�����V�*���ۙ��$���������Y��bI9?��(V��E���E�����d��ĎtA��J&����M��Ӵ��93��A� N��1A��/%�������Eڍ��L$�z�'��%l��f(*�v\����`Ŋ�#�~p����s��\)h{��@;w� 6>����/x��k׮��i'��D�F x�8e��7�#�|ۙnͤ�o)s�uԠ[
}fѝ�e�.|�\<]�lYJ�� �-�,[;ǐ�>����ݻw_z�o��Ğ�{B�a���~:}�ӟ�M��Sz:σx�\O"��G Åbε7F�8"�U�/�{��m��ր� �����)��L�T!o�|�2Z�j� �{~{�4p�<+d{�u1�?C���VOryM?�2}[����3�/h�!�`U���Jؔ�R��@�A�FW�ΨYҪh�[̦,!��pTq�f��"3�EQS�"�1]Ӕ�L:0��P1_�2�}�	ͨ�G�� E�vwj�[��D�ڄ���g��YǺ� �Z�&��Άǧ����N瞻�����B���
�:tr��0����~<����W�E��\{o���7���i�V�xO^�[�0��o���ַ������D�k_���~��_����H�1E�Px���a��^A<�# �A�Q��i�������F���_����+�2+[Q�dp �U�V&��J���s��X����ɀ�O:7�ھ�dՔ���B���!�Vڡ.�W8�V��+��N� ���<89��oӯ~���&&'Z�[(���w��>򑏈X>0l<W<c����8�.�p6|tP�@�@FT)V��_$�c]��O�il۶m۶���N�jl�jl��m����'�Y�g�]���~Ln�Ά����.3͂��02^ �E��hw�e7�w�6�`��}U��St�1Bҍ�ڵa�#�/��N=�J9�Uk�0ٻ��e|Zg���?w�.��e;�#������0�NhE&w�Q^�+��
�E��
p,�xdqQ1�Oy,W��D�%�l��5�����vW��`�R<����&l���«�X�T��Z	�J[��q�7J��Q�?��ozt��|�T�_�s��h�n�.ێ�zsU�8����yӓ�\��\��:�v8=�G�)�����qW�t���	F�
ӕ�ոSxܝ?B9�m}�߈`<y�9Gl��~4A�Zմ~-ArΣ�'��9i�cC���)f������o��'h�Te���K��h3'�Ge��Atf6Ia6�%W!�/��jP�.;7�:J%�W��(�&��O<�����Ը08�N��頱�4��f�kEף�̷>my�n:��mo�~)�o.��e�����ҥf������ZI�"F��R�I���o࠻�;G�}lع�݉�Vn����@-X# ���� d��������+���t���|�E�|��uL��	<.��O �	��:]�n+�[�}h�ɷ�K�ak.����D��@٤�Iɟ=Y6����9'Yʅ�ҐL$z�p3�i4|/�i�~�p�S\��K���&���&��O���[�W�'�Վi$�MUVWz��.#��|ND$D�h p�A:��2u�ۉ��e��f_�ڬ�c{&`N��e��ή�Q��}=��`,7Kl�o:OT]�m{o�1�A���/�^�����kqD���7V�P���i�RO��!�Yr�)�2�Eh�%�.��$�З�v�x�������7қ��;4|�1�cb�\˒A�uq�PX�����k��CTo�B��T,�e,�A��'�>�K�������&=�`��F��Ӟ2!�drly�w0�:qs��{4���;A��N[�&�����mj��8-���<!i�.��C�PP*���K׈��S98�X�݄J\�!���2����d$�Ǎ��\Pb��:-j�'d-M��i�����J*��9�V]F-�� :��o�飍קؿ�����	�׆1�����F,��u��Ə;јm�����wu�pYD{`�����GQ��#�?���M���������Piz��
=ej+� �_��7�}�uyM@�R&�O��#agd�������9Q�����~���[l��os� L\LDXeee�~w�
x���s��vF�>6�rW�W���2�$.i�]�)�֫8W����l�3��!	f�W��Z�"�1��l��������t����dMmM�Ɍ�S���)fa}���%b�g���3��G����;��&h�8+�R�g�Lؼmy׃,F����f�CufL�����-�:|�=ܽ/1�.��$B����f壊�ߌk����'Z1H��tc1����\�K��ɸ�J���y�d�u���SwP����).�7>.`iy���2 �s���1��k�y�W�����+�ێ��z����oqK�q����o�5�/��4ጶ��x����{+��lQՏ^t<�&�8dv����33�G�#�X�@B�T��yv68t�4~��+4ߟG��Jo�M.�� ���?]�����}6g��3�P0�n����`���w]eD+|4P�4�wR� ���d��{��07�Lc
�S����U�&ϚUT��N�@�*HifZ	��A�$c1hI�N3q)o� X��Zi;t((��v|�o�:�u��Sz���O�%b��y')<���/�˹�K���9���ժ�o�ߴ�r�>�&#`MU/D
P� vB�Yj�+��
n�b�"�c� l�(	)h�������	l4��w���Dq�<�5:x����;ČH�m�.����3��
��~����4�MC��]�=�x�ߌXY+�ۧ���\��ӷ�5��J�'��kR��G�4�X��I���8J���\��Y���8�t�z�������?�)�l�}��1#�
�{��}޶�~��B��I�
��|R]�__.�������p03����I���J;4�w���E�����^+�����i�2�~B�1'�ZquKgc�:���采����g_H���~9~>d��ep9��²���ez�/���r�����TǾm(]� 5���V��O��M����_d�q�oLo�<i�C�;��q�7x��o:�����đef���E�ZYυ�;�k�Tң��g�V�_g ����ep��fn��� �&���±.������/��{{�bF�� ��zJ��w�zخe��]Wn9C���vo���+L`������Yx���,�*^�6*�xpI���b�LU�oWe�0�w��}�B�պ����c6��7�rCgB�i�w�������M���UI��\z!&ŢЉ��S��8�>�v׃.�Pp;���t+$!.\o�˅mx{{��
�:~����j���ͯ���O"���r�����!��X@�D5u��Zݝ��;���d�~��O}b���:"����`�lܜ_��列�B�����[��N�J)��B(M��J3���G�?�f���XT��|I���[�f@^,���Y<�>,�7?]g_��=��W�:?U��m�.����<��g�fij�՝�¬�3�Rcl���'L[�h;�8ݕ�/
��:�5Rƺ��)�("��`�K`f�H�I��BO[hhP<<]��y?�����l?�,���e�>��[���IYG��B�(6s�k�C�� �j��h����@>��q��o=��$)ߧQ=a�����{����2_<zu�!YEu�\�׷�̃d3pٖ�a�F�D����j����p[z�����͘>4X�{��	=�iD5�ò��Je\-���_�q���8�y���c��:��a���Kj>r�䦽���� n~퀹�"�+�����Wk�-��L�ٿ5>j��b���U*~�ڥ�T���UU�$�gW�FԻ�K��h�
�o{h�C{f�����d򳙡���� zY@E}F�[ei���	dl�:;ߝ�䉽 �/�w�Z�ū//��g�B�mmy�l��d�Z��JU�>x�x�YM+Jd���̏~Ne��g.Ԍ��ǖg����xH���_ME�ʖD�c�X�XlMM��%�"���U�����@ �EF'�`K�4��"��1(5>|�~������L��k9��7WY��)��/���s#����|r�;m�0V���b��|,j�\ۤx)yi�F�my�KJ+u�Q}���=Uӟ0vz�ʁ$Ў�!��*(������U�DZYg�x<S��
>+�������N)�ņFZH��D$�M�vs�Ǔ��Ǒ�g�u��;̴��W���ɬA~���}��O`�W��]�9�H'�[�M�u%Xa�`�Ji�b!��z�ʔ�b�Y�Dq�Q.g�r4�Kt.F��y���S�WWXV����D%?a!��zzK���`RW���Ɇ��J[gs�?["[�N���)(�6�����U�<v]�j�)�lwL����� �r�*)�u�,����O�ϳ�0����N$8s�g����\�0���x䓠�����Q������h�^���y���G��$����׏�wn$� �!�E`
@mpUHG���M| x�~���$H�&p�'NI���+2޴��j�1�=�pAqRG�3�D�]�>�М��EU{���{t?�y=@i�{�ؼ\l�9���V��zq	�;�����϶�3��h��h���M��>њ�9q�v�Z}MhZ��V�ځ����769lw��DG�*��D�ʠ3�q1����8�a"A|�}t5�6�%�Ub���� ��#~�v}�x�	2�=���� �EBR�Y��O3l�2'��J��(G�96}P�>��P�N�a����vVW�#N�0�c|�����(�x
1[sz8��7�?�Xp&Z���b��D�r���5�)�
�^���C��̱n����NJ��~�m��by�<ff�v���� 4,�����Bp � ��)���\g@N��gV
9|X��l�j%o\������!oM���R)��T*��ʝ�bVݽ���s�۶���1���S��t[���?���E��z�j�O��5
.��ڙ�N���$(�G�������m6X(�!�y*��r�����M�B |�+��;�f&�ٽwk�dNqf����=�|��U�ج
�5U���@���y5[s�����D���).	�������E��R3ֺYZ��q3,���
x���4��w����b����e���:bh��{.$Pi����*��ZX�32�
���)T�ݬ�=	�pIHf��P�0^�o��~5���}��8����5i�e��{��S!F����"��*��b!>)��eQ�i��d1���N���z�Ԃ��p�Ȱ�̻��X.���}o]o�blf��saM��]�>tڢ�N��1H>;`�$JA���/~��?���)�Av����f����6e�������ʁt ��U�� F�0(D]>&�t�[���#���*�6a)3?au;F�1Ra'��r�!�m�����<� G��K@18x/}}�f�^�5�Ū?��꩟L��9|�S�M�6��BGMK_9U��8~�<�S�C��������sd��J�S4�9��q��f}:��h��mF
�|��f9ҏ���D�� ���k;q��	�lKV���Ĕ��u�}�Y(|��m�����h�p<�^�1�&��K��m����7��F�_�������on��uėN|Y~�p窪q��vF�ϯ���D�-��R���[.�~�R�_r�n�}���.S\SG;}Aײ&�#nԥ�P�����`׿͜�f+]���288����J���Gk�æ��Y5�,�K�=US��ڲ^��|(3'1�����1:�ㆈ�p���m���*j��Ż�Eޏ����d]�4��e���,����T)�pP����㥚ŏ�3�g���M#�*��劮�"��sҐ�=��O��;�QT�����C��m�	��%X�m�^��g�ץ	��Q��_�.}�����,$���݆m����}�"Y��5��������=��6�S[���v��oP)r-����y������i^�&.�w��n��GZ���n�Q$9oV����R�sۨ�=�s��3�:,�-M���c��UW,K\�m+l�m=�l�Mytu�N켙e��"_�k��
��ɵհ�7�(�y�&3��b�i)h芩�mnC�-�u*i4!�-q��������K�W1+�};0$����	zO�_���Kׇ�1y������6�T4fv��e��G��/��dT�U��(�yz	�Ȑ(Z8��oA{/��&Daa�)�NΏ�1fM��*�ʆ:H���s@^7J�t-J�׊�Q���C����X8;G'�n�8�9�n`g´,4.&=��R�ʄ1���<�>��7Y9��uɤ؟��)Q\6YɄJ	L׹�5�\n��Y53j^�F��3��O��.�_�a]�D�pu��r��c�͸��>��o��>S��[�:-��4�E ~�?����������-J��J��Iɸ�u�.C2�yt���1�w��a-&�"�������^���<[7���� [������ұ⟸c�ɛn��G�ý6O��HH� �1�{��J�W�Hb�q�AS��
	�H�������0-����i�eד���]�B�zU����rf2,�:�u��-W>'�%iX3btD�|��;?_�R�@�� ^x�P�yU��{A:�/�A3����ew!� ~�mi~:���,�2���6a�����@�S�`M;˖���F�Fk���D��V����j��m��w��WU\q��H�az�t���C���`d@�×�Z�7���M�����<����9�2uN� ��sU/=9�9Ӯf�%/jE5r��b�����r=a��T�#���'f��e�PH��_�\�:M6ݕ���H�f`����٣��`��m�,�n��9������ eÀ-��
�����3�d�ρ�I�M�	���i��S��Y��ף��A3���{
�8�xw�z0Uo�^{���<"|0+������H�$A.s�h�Q2���-+�P�3��Ue���B0�E|W�$"pU�K�u^�E�nV�M=�h��//���U1�������Q�4��um�XCk`��߉J�sa�`��J�sѵIW��|���O�B��e�h�]lȜ\�X��j�42����Aq �m)��H��U��B+,,T5�is��^ks�ȑYs�|i|�lX`�N�x`�g�(g?�-�DrA���;�E8�˜ʃ"��9LNq���΢uR�Bm̵y�b��z���3[�$B)�������o���O���˩`��d6����L�=(�N�j&Q�`x�k\I[҃�ښW:r&h�
P?�XW�G�7�H���cV�����2>� r��];���ol��ᔸ����d�d��E�k�e&�o�ܽ�I�>�x��:S��/u�=����)�)�0:#A�>D?�斉��7�����v��Ƭl��k�KF� Hrnّl�j�@�`m�
h�����mڡL�h��)��f�xS�W��j�P�?������v���CM��-��<��L��X�ĕ;0��$ZcFA�s����v)��Y@���L�7�Ն�B2�q�@+��JF@� N���3-WZT����������Ǽ5�����\��?**W���?)��f�NV���xo����^}�n��#��e��J�O�����I�S����4v
C)�(@�2��,�����h����@|3a�#!����Ğ��/���嚷vS���:�"Of2�o����3͗0E���s'"N��6` ������t���� 5fR��?P]�t�p%�p�$o�E״�c��$���1���5��'l�f�ަ|[��a�q�]�K`�	)m�:YT�X9�L^3z�AJؖ¨�h	����|��:m_����үdm����G,~�g�ZM����~��ʊb��\bO��`�	A��Lx�+����������b��)���D���Vx���#܁nR`o�_h}�UZ̠��z
D4C`,CO�!h����}G!�T�--S��
�w�nu
�L74w�s��q+�w�dZ���0����N^�I>��_��{?#�:��&�2���5ui�~MT阖�-Q+��;�E?Sf��a��
~�0�m�;hf�I/� f�.���R��\FCh��"8���|� �Dp�ZU#�n�6gl�z9�Le%��G�Ϙ7�^M{�C3r�T�V�89c>u�H{�=T�����d;�=��s8�k��~.�[�4��n]>(H�?�U�HYJ��/x��G}#�nT�X���C�@��Uy`Z�#��A���6x�i����%��͋
�Eu��퍔5�r����i�r��k��f����f��Y 3+/i�0`��U;r���N�G���� z"�$ ������c�V<I��z ��e�S\S�
pu�61�i�����x^�BÛ\~�s�!���O$�߱�P���/����B��V�M��^P�Ty7 �]�+��$�c�Ѵ_;��J�B��.�Ʊ�oX���d���K](��ׁ$І�v�g�J�"�&f ���ޅo�2�����4�8������)���=E~�a�mO\'����5�q�*Yx��w�	N�u��L�tv�5gu��*���\����/a d��C��g��l���G�!���zn/heAM�B4\��R����d	'�Z|�
�ndd�*]z�A�7F�t��}>.v����xr���E���N����3HǕ���w[��O`?�$�ޛxV8�sۖ���R3۷{�Rd�q���xH8�)2�т2�0���2^#V,���J�S26����TSJ;��oz��we\.�C
 =�!�ʫ����V߿A�Я�hk ��pk��*0s���::���;���.������Wɜ��x_���w]���0��(�G����FՉ,�֡�;18
��
�
�ũ��Gp����T�u��j;zc,�D�.���������)���ڵ��S�Y���߷��2�����{��%��_�Dlb�ߝ����S6\�{C�e�Fh�A��a�` \=@����S۱���Zl�
�L�m	���\��Z��=�=|,TH�̻~v�q;�ƽ%��Ő�Ri���o�_@e:(�BB��/�:\]�-x� ����Pq����@�Q����|xO���ܩK�L=����(,h
����d=��g�!=�Ke��>���I��K��um�D�����za�r4l�ֻ4MK4�]�.�Կ	e���c�gH��f?P<�Pͤ��IU0�aNS=d�$��W���^�&�����Oʋ�6f9�D���-�U-J6�1���Y5�.Yȇ��V66�����a��=N�2f�
��n�t��z���io�k��?}X�:��, �|]|ʌl|l��7��}6���<�P��#��~q/xf_:`M(���'�$�GI&�d�����e��K $��?�|�=�T-y�K�.G�=Ii_�k'����J�S�K�@@V����t����&�AνO d�c[wVKLm���>p;��s%��h�^��<{�Riu��qlCT��ǰI��P��~R���m�5�Zw(�e,Ў8�[�$�dq�N��VNL
�������������S�MN����4]S����"0 �źբZ��.,ڗ�J'UڦN���Ǘ�[RoO�Ec7J�)���55�]	ژ��3���z.1@}L%CE>�gƘ�X�+�0#*ϓ��F�Mj�0��ݰ���m	���[^O��Ŕ���V���:KT�3��� ���ׁw�o[��?M�@��,ߨwa���J՟���m+6J���a٨2N#k�@�=�SK��=�r>�Ë́aa��p�v�Z#�<k�"gU�)1�����	(�0���w�[yz�}:~��u0ac���76:�9����MN*`Մ���.6霖�AQ��\z�)
G�1�	��	��+-g3��P�BT��D/�b*�J�B2�Kr-F�s��D��,�G�خ�;��"<%S�I��R��@	{((J��A��O]\� ���
��.��*�U� y�L�*Cm�5:�س� ��/N���xS'`10B�)1�\�N�l��Y8���S��Z� z���K��{��z��h@��Mk���O�\�Ј�&��Fb�9��v����g�"B�A���+�!�",~�����~2q)T�>�@�0׻}�B�I��o�y92�A�!Q���, @�+���Q��	L�I�i���7Ϟ<
�z�9tۆV�M���l�0K�����ߡp:cr�������UBQ�.n�p�(��˃'o�@v$o.�w�j�wk�o��x��U�+z/��F�\�^�]����-M��ad?C";�A�ʙ�F%� ;�L�nT:`ن^;替��14ؚ��s8� �ޜ��g���8��~?�UbD�Ly\EB��J�%jN
_p�����ToC���^,�����_j�kK��0���.��>8��-�E��"f��KM���� 2�L�X��p�'V򺟕������多2���"���Ӧ{Q��n�U�n���ND��Q��2��a���%�;|�JP�X��u����Ep�u�rh���)�>����i�$$�u��ϡ�md�i�roXև�*;jZ��{�N�~gQ;�2j:�k�}��T�K7�i��"�����ej����~L��4:���!�
;L"i���irX��ha6�h�!�U�l��8����1X�~���*Dَ*26�@?���K�B�j�~��=�tG{)�Y\]����K8�%}�N	�0�=��>@%(�������
@���J�ڣ�`�嶅Y
)��=
��l����J�i*k�.��T�?%�,e]�K��'��Td"��![Z��P|J��5�51X t�L 6�O�4��%��.A�n[t�}Wp�g4�$d#T1!�L�����&Ajw�t�V���)K��(A 2�F,`X�os��0��/m�Z��(�2k(���,�VZz�U��-(���63{�$�/�&=��+��gT<����J1�9_xN�?���pGl�+?a�T����c{%$OJS4-�g���_�U�M��,��V$���c=��͘xmi�\�|�����h}�أ�/���(����)h�����Q2��M8}Vo&�|w�,��5�<}�'N���6B�BV�/~������&8�9}
:�Ya�.bڤ9�3�!Z���X��ݓ9��Wf��8�w����/N�H���	>Aϙܹ�s(���@J�CuAONg7tұrzꍃ��!S4b2�㿽�����E��-������5:|�cgc����|Y=u�[E�OR�)�ϐNпF%2�Z��C�0��� �+0i�����ꗩo�٤��TP�E�Ƹ�9���_~[�g!{�3�SL@��Ѳ&�T0�Ӌ�cݛ^�A�UؒXSƃ>~=���sw5�@v�
�C?��V3���{�.T���1�I�g�eNGz��DїX�ٰ��&梢t���θ-�IX���?����?,�f��H��Q
���>N�A���k�M�ӓ�~:/��Τ���][+��C��	������ɞM�l���l:M��EN]6��x��k��%�i=�t�ەB�r��&p���y��(��)5ME�6���S��aPf�6{?I��ѱ�ߍ���t�>��P#i�����p���S_�'���*�N���;O_Bԝv�z�~�g���ou��qq��cIѫ����x\��E��b��8?� � G��qꙆ�"u�te F$~�� 2ǀ�ۯ����+tfr��y�;�k|Y0ğ�`'����j+ܓjA����8��G����jr�,�K��nu8��vk��FH[_ 2X1��Ϡ�;�/1�,�H���5m˻C���_�]PYznM�=�\�\�	��s`00r�ET���o�袭)Q+p��Ǿ]��g������Oj�m[6�s����������'>�+>���Q1��YJ���{ztδ(�Y
B�F�?�&���ìF���t�qJ<q��&��b!\����	����t��Gك/�7o�Ơb)|xDx�.:�ގd�[��P0�#���1�4�_]�{+����u�6���?IJ>@BZo��">��t���V�ShO�>w�zv^�֛����߻ww�^x�y��Ձ�y���?�C�_��fR��#cy.�ۏr:��
�S��tZ`n��5�,�k{�pG�r:��+�8K2�E�B�&\��l?mzװ6�"d�لEDH���@���8�1h~h
�����xGf:����GȐ ��o��C�N
�*L�/��?١������N�m��\nV�����Ǥpm���P�R�ߋ�<G�{�v��Mjo�U����n��Mp��x5goeqQѻ�B�tkM<m��:��b�����KA#��OK�m����#��>^��iO���~�=����p*}>6&l�y���p�v�;?>�{�~�c�u�������ܓ�����8/���A���3A���r�P#�j���nme�P�t���N��HX��ֆ����C�|���8n�|_a�k���0��ɏ�B���F�ؐ
Z#��Ke��Kg%ܫ��z���V#V:V&uzv�hy�l���OY��y�$�/w7���a������Ko*&��6Vnn�m�Q�b����9��,i;��ƛ��b`������a[�.��&��[� ��I�TB�R�B'^Yl/w%�͍ B��2�1�F v�D�ߏڵ�,f�O���������	�s�?�΁��v9Lc�-�͑;c}s�.���w7m���N�'�+�" ��*{|�P���@ip�c���빹EEA��⯅��JD�+S�x�`��K��t�eRh��#�?����?�"q� ���� ���?�%R���!-|�!�S�S�f^�hͰ~��D��ֱ���E82.��}ѭ#\ӈ�P��+�r�
��q,��#�B�\rE�
���x�R�eN>^���s�zQ�G���z�e�V�L����x���3'�$�ߍ^�R�I9�y�:��e��_�.��p.�6r��.|����Y���2�[��"��w��'�T�aHꚛ�ۆt�K\��:Ĺ�/6�F8�J��?�w�[t]�-��*H:�M�xĆ�-se�\�ҶoAg�Q�{o�9g0�R`��~��Y/���e���T�@\�IOحL�:� �zv��W��0~�FT�Ͻm}�{}�1���w�ގQ�XXP���x@��а�%K+e�f������G|2#��kl
~ݎ)�x����`zʽ1�	u}���60�=��]Vӏ�<MƦ1�|�_G��y%�C�a�;)�m�yS��.��*�����6yFm۷�<G���P�ɵ�-�q�`?>>��	��Rʎ---���FnP�pџI�?�_��/%��uu��0�d�м2��v�%s�3����s��A;�Q�!<Q�W�Ģ����u\�[8��u(įlK�~��S�X?UJ5�P��C�����K�& �wׇ��uIWN��pZ��������לu�t��S�O��Ch#x�_")��8�H%��Z���xv�H֑I���1��>�9@x�y�/�����ͯu;�N��g|JC�Qv�� �i�L�-d��I���y������̬~Y�8�~�:����Ѻ���]�k�V�i|���Eg8OI!?=�a��&�	�d��(��o¸���^��n�+�h~n��m�~ܑ�W�wO����ӶКS���\�+�f�Gu�B��.��t�&X�OkR�+�L7�/jJ|>�=��ن,bΧ�"�״?��0'��>���m��4鉬a��=_�1^?�÷�z>���4�b�0��R{�hjZ�}��Z?6D��oIӓ5�y��B�)Ψ���(�	�k�O���I&����p���0�����v����p�VvÞ�2�x+9�Bd_�o%%��e��ջ���LNٵ���h�7}b�If?i�f/VG<��p���Έ"�\>�k7�X3�]�Ӎ.m9kA��ȥۯ�C�^�Y��{h�7l�,�����X<�\�d70}:=�uOpIZ4qMT��J��������K�*g�����Ւ��C�_�o՟8���a�_���`�EKU{U�|�x�L�Fs����:���90�܇	�#q���bM/ű��~�:#��ӟ�7N[V�I��r? �;��Y�/U�/t#K��(4֓I�"hf�k�jFky��|�����﫰�][ɍ�EN���k��d1�:z|����w�g7�<� �OE���5ٷ��*W��F�T+����d^�/k�H��l0e��A��1��E�
���$ [�y�����F���i�"�>�$  ��Q�X�Û��a-�^;�g��2\%E��㫽���>	�+#�>���ήo�x�~�K0����GP�(���e;�Sݧp�$g��~����T��Zϱ�9�����Z1S�C�['39��B��C��^�ޫP��J�� L+5����O0o�+L�/8wQ�?'dT�C;�q��1�f}ҕ�t�/~P�Xؽ�����Q!Vu5���@ۿ�bL�8~l�<m6>�6%�:�Cť���y:F����hbUo�b|o��~-� �މ]w(���P���G���t�K3�x0�YZ�"o���z;�B� [���e�Ŋ����ð�V������_볠$1�wO�l�cgggp�A0�f���tx�$Z��#�7z!�{Oq��-�_�dzi�u�(p�t�8p��ly�@��|��y�O�%	�����p�� �B���a��~=�H��''����?|��CWUI�@Tb��)�frXn;ʑ����j���v�����5�o]ʹ�-��C�r���t&|���@y�v,-{��6%�ƃ������ )��Ugu ��3��|#���x42�c�j�a�o���j�W9�r��nv��Ɓ�ςR�ظK����멋����Ȃ��e�j� ʂ�^�޳$j�:����i����~Z���Z'�ۥ��#���}H0f[�Hƛ���;�^��q���ý�����L㧘tjo_@H����Ν�������J���-H�$aJ�-x���������$Sq���������)X�`E��B��|��3���+�/��e��Q�8���%�C���a�/�~Y� ��|�б�O�Q��Cd���\v��}DQG�U�|�Qi'�{5L����N�P�XV�>QP$JM5�?dI�m��%qs�-h�|�r]Lր����qvW�l1�0p���C������Ye�o�"��ݶ<�|oy�#� �AȇCG��&�X���r??��]T-'�����2e�k{·f�+ҡ��硾|0�;���?\�w	m���1�B�p��t�%TPA#�cC�o"�n↛B%��)q��K�/�R�}Nd���K)�j�`�4H��i5�S"b�i�( S{�Ar�F�RO�gyC���V��jT�=�"������3�|	v�$^_Z
|�ȿ�=3�y�Fam���AW����~|�!u:H��DU<2^V��J���D�����t��T�����V���T����SY�*V%��$+X b<��~��Q��r���%X:���}ٞ�Nk e�T���A��Ǉp�����Jx�Y�x��@��׶G�UZ�9�����6��z䭜���D�,$P�oؠ��+�y7��~n���+���;�8�kT�:���7�qP�}����/`	��|�z�z�4��H)%e�I\Zb��&U�D�7'�r��e�aŦBMs��1�#�)� D�Δ�����g��yL����I�,��h��f�F4��rY���R>�ҽ9	PK~_�8���Ԛ?/9�P��2Խ�֏�*L#転�)S� j��SE{yYP�#3�v��T��c���ţV���c@��"ҥ[�hp֚3�j�����͞�Sx�	�d���6�-U��2M�>�L��Z�M���'Bs�+*?�28:��nT
��mM{�����\Z�g�cȢ�W#�^�&w����f�oV`�iY_F��D��o�yˏ����]���֙1���a��57�� hU".��<-��������	��o���5q�q��W+�q���tZ�i���b��`��F���?p���=*V����F?��������x�a�	��4z���P౤"X�%U�x$��9�P�A�e�z��Ή�|��٩��"|��-=t��2��[[�Lr1�p���<���^B����m�ظڶ4�= ����[H)S���hhj���%׸�*6�iϓ=������6��k�[5�5�`��<Z��jW��0�o�7薝C����B��6E[���5M%�߀ΐ_Qk �t>�x�ÿt>_����8\7eM�Pj���#����BC�#2=���\i���;X:Cm�pG�!',���횐%G��g���\�oFd�f�Z���_�<98�_OJ{�z�~�
��O~\�T)O�P]��NK�� @�
�C	�0�Z�F���#WCG8Z���j<�䶿�f�3�ܞ.|����&���� '��C�B�oB�	B�P.aNT�6�ߠ�Q[���8������pH���4�6�T]on���ĘQ�eq�W���jP�+l����] ��a�NO�z%�9��F,�>a�Fx��8�]���������(��eݴ����##���V�M�}~���%^�H���T$jh�kG�����[V��st{�͂��S�&As�"p����	=;�����.�\-�KV��I ���`@F�ۂI��A� "ZS� m���euJ�?������ܠ�Q�^���.\�(�Ǔ+������.�>^��`'k�Y��v3�\N����?�p5#����!�:��`r�涐Y"S�¢�ciw��z>�{"�1z�ŀ��A�;f�aY������qo9;���P�h���E$clS"���������j�ڥs�7*t]��t<7��h$��"�:����&�FX�u�}8�i9�O� 'c�բ��2������v��p�����1;�%���&lC�f����������>��6��֑�T�'��?W'�_W=�~7���-���h��	�4Npwww�ww'8www��ݡq�hpN������U�j�c�U��]8*��2���x.q��Yh�K�.���c�0ʭ7���}�"�F��x�a�y���q���}Zܧ���ҀP���gf�^���V�K�R�sٗ���R�g�V1����w���	��f�b��1쒐g�eu�@�?�&+Op&by���x}9t}Ȍ��6@j��CYݲoݒ���\��~pE������`�c��u��[�/��W'B�~�9|�`lp;����B���58g�%u:��:��6��dX�c���%�o�d��{�$s��g��?�&��H���sV���R�Q�܈(�+��ɶ�㳛�e���B
,"���>��wf��fo�v������3�5h�e�z��e�L1�L��y\����O��W�<�I4Z.J������p��r����*%�(����S8��7e��PE)�������KЅW��	�)�����v�^B?��N�O�PzF�;�Xr��n��[�@-�פ�L2�U��?�T�>	G�o�Wxq��50�i��ֿ���Y����P$j*�]�0�W����_�ߙ?����C��ŴPqD��p��eF�O���]b;��s?���B�ˏ4�YZ:~�X�7T�Id ڃ��D�g9��W=�2u�!��;]9S��=�;��&d����4 +XJo�zzm�h�����`��}��ܞ2!n�{�>�̿?c��LL�W	��f����T�fU�u���f������h@�������킝�/��:�"K9v�	���dB�C����'��,�ڢ��X�p��PY�q�v�K؝Gz5Z���s�S�&6��v�d4��i|a�����Sq�<����%]�s����3O@f?���Jm�~��w��q��/����ppx��c$����~��yk�f> 8���~��)1�6�)��A<�h�v\ۊ����ӈM���8����yRd�&V ��������
�6!˚0
ݥDt�D�g������<�1j]��^��B���Z�Z.Mf���l)��R� "c�D'S
������%v�k /`���Z�&��`��i������N����Q��O�����]X�#�g�qɯ����b34gk�!�g&��B���qH"gQ�.���
���,ҁH�8�DL�RX�O�h~J��s�z�~� ��	����gZ���Z�.f�tԕ�.��U���?��#���¨0в�2�ܖ&	��������Ls��Q�S���%�<;��s�!���-�r+|Y ��S�~ڱ�Ќ�ݡ/�#e�����kH�S4�-�c��d�.���.��Z���0I[��x�>F&���9����Wj̖��\(-�&[�d�@�ϻ��~��F����W)��P��s���b�!�';:�O�`u�	�\�eiE��n�� �5� ���*�̼�HM���1��p/0R��,��1�~O&ͮ�~W���==.�(����^��� �J$ ޚX?&�)2��n^������<�	1>���Atч*z�v6!��3�I����NK�(�1�W��B�Ai����.w���;��˶z�'�4.��;�ҽ<쟤�?:���־��#��Ϣ�O'�Иgp�9VzQ�@��훀�I1D����(��@����*$�
8k����=��鼦5�е}�d4Μ��#�m&.v���&���wU�iF����
 ��Os���گL��nk�1�B1
�����T��<L/��^��q�Y1-Ͱ��9�|=D����O��
ZKX���R���_���:vն��7�[jM�Ͼ�0}^H>��6����]V��JE~����6�A���zm���9����;�� ���N��!2֔\�)N�0�W%�$T��j��)2�^�88������!b䂀jnN��۸���h��jt=��8$������ͬ���!�#̌n|�1!GO�s/7����({��
F��a�����<=?b	�+q6�Ƹ�%��+��=׋H}l>l�Z b��ޛ���e)�~d�)]�"N࣌��Vw�E%�kvW����-��~�̈́%��DgY�B���D�M?��zAd0q-H�g�=��K����EV��=Pif��s��*ǆ��Kd�b%u�µ���i?I	��6��Y�L�I+?<�������>_K���������dP��M��'(�H�'�d5e�)#_;���-'BE�8�����24Y�*s�,��Nf�ϓ��w?��j8�t�y��P�s˝Z�c���� �T��6k��8~U�s+��32���O�v�g�[���Mֈ��H�9q�a�[�-��&����.�� ���7���.����6)����Ď�|�h�l=�Z�Ӟ��hH���>�d�����i�� g���7�~.-r������� � �5BoH[ o$��1��f��q�6p3*�v��s]�%؝�⼶Ѽ��.I��x��!��^����ˤ� �>La	�U�>��sfcC���HF�&��e�{�ZA��HQxX�l���IU�w��I#��=��7�l�]ѣ��s�?�b��&�_G&�����s�=9�|���)ͅ*�Y�-,>�����o��*��O�GE����c�?K�K@p��Nɟ����X"	��Q)�������h�S��$�7C����3<��k�B�n����ꗫ��+=����%��w��/�];I�qZ�,�����gI�Sh��CnyZ�Í�GdTՐ�D{F��o�7�jf�̫�2�����P=�x��u�z��Α�����~�)!�R7��x6�Hq�7�;V��|�YȮQBצ&��ä��ޏ�^
m�Ӆ�T���a����l��1�I�:�x��m�����tˮ���c�4"�kC˫e��4�GN��>�wy��n#���g�{�Ƈ�dd�[ˊŜ����t,`��c�/Swՠ�+��44�~������5	�D]	kÏ����Ԁ'���R�����S�8��o��mGi�f���/s⨩G�@b m�!�)2͙�d0��n��t��p���(�V*<�P��ڂd��t�(��O��]��e����p3� ������ް3� ��S@ ��g�t�J��a�j
DW�jf�N�G��Eݡ�����}wf�FC�0@M��[��W��N��Ƃ]��.�P�����ɺ'�j�:t~������#�m����3���+:�X�ŋs̛8�e�z�Y����j��=����'Z��dI�N�����%�Gs��� �=�F0��2�5�c].�2���?"�8�9�g������D�{�C�(��[i�s��d[��z��yJ���\wRJO�G]�p/�n
u��_mK^
�x-�L��=�ѝ�;��.y���WE�ڌ_$���ݥ��"�I{�ӷ55i�Px<C?"����o�Wu;=.�������r�j�V'NM�f,��n�K#�GC8��2m	<}��u�/X� i���b�c��g% �����F^��C� ����w�|q���	5��[s�B�`|��ɯ�W���x;,�mu%^MR<��q :`�`G��Q_W�U��w;�o|�zD�|�7��
�
��=��۴�.b5�r� �M���Z�J�5�r!���;}ӆ'5�W����^W_�SO$�(	 �`�*��\L�%���PN�\�x�>wM'x�U���/,rV/�#4�o��P0^,��y�hk�_�����I`���?����[!>��|�w�o�Ib�}Z���K@��o�#j�,P&���et1����s�����g����N�J���ޑ�O����ڲ�"j��X��wh7����A���TƊ;G��5h��`���
�H!A��'<�f����bJ��˳i�	��R�-�o
~���z��5�#o���6!���5��F�${5���v���|K��J�rK$��By���
��]l���mQ��a� ȃ��|�h�<4�zk���'�c�M�e�k���Z�����|�~˚��N'�����@��SΦ�fkvSK�)v������\B�'_;�e��$��	�ވ�YۖVյ=�7s��(�;���"�
]�;��}�7��9{s�/�@�{�D��t��>>>F���¿X����?���m?�{.++��H���@� �~�K6�f�"�?t78xQ��岼�����Snz,�h���?go�|bH�Z�a�B{p��)����ŗ��U�!�����U�k7jZ20L�h�~�g	H�Կ��f�Jc�f���3���d]��i���ge��
�e��Y�J��O ���qP�n@�!D"��3���W�B�N4Uɼ����ظx�+��lEE��yI:���k�~���zD���t%����߳|�UW�[;{�[���qn�ѣ�Iuc *�xol-���:���;���s�׼����2"q5*��t� b(6���6��^?�=�@?�-D�f{;�]5z{P�b �+\��أ>��۹���4�<M�`#�ne7d%����DP*�P�хq��8{48tbo#��������'�������>t�J�Y|�-�]�v��/�ױ2U�0۸(\���1�y�7��tO%�O��](�"�`u-4��H�@hh��^e����t�?\��ro�_I"����R��d+L�����}M�L��O�%������PE$2��y�.�l��D;4����E0��n<&�O��E��z�=xx2�G[�&AB�;z��:��������Q��Ɲ=�ԋ@+�*R	�ǂ�>����S~��q��i��I�"��L�r���"ڼ����?#`#�����~	j鱝�ݺ�5�ĥh�j���U�m����Z�+�G�ȣI�CZ�>�&�(����(���`��`��Bv��DA|-(m/�Cs���i��C�QIMRa�sw/_�������0�|���5N��>�$�Q{���1������w���D� 7��FU#�]�v--���޵ez:7g*%?��SK�TA��{�ӉIf�$%��x��,D_��8V5�󰍌h?��0������Ϫ(�����Agc�뷡����� Ɇӄl:��ϵ�Qʁ�w�F��bBo 0g2t��ıo����q6^�',����#8Y�y/&�y�t�9�aN�[������@´nӁ��>��`qisfG�����η0zIe��(��=�9f�8D���r#iw��AL�fJ{Yb6�-���s+L��j�!��#��]��]N��u[�޽u{��.GJ2�Z(YC==��z�ʏ��L��/�gY�q��t��9K-�q���e Cuk�'�#a����>���">qq�N�zOgqbL�K�,.�pWh�U�����خzD&@�9���VP<3�S�ڒ�Z�J�u��,*����� �ʍ6kң�'����6��U���ހ��x���{��<ط�2TƊ��VCa�1���n��ˠ׵f�t�h��t?�Xwz���0_��
f���͞���h�x'�|Jup@ĕKi�.��y��5D��W�Q�%����e2
v��Lb���Jz�L���_'�J��_�� �(�"!`�XQb�G�k�kN��ф�f��I	?띡�N!���w�y��9�DU��!�]�I1��g��$�>TCt9Rф�Jlא��j"�qu������jSέF�.�+<��0N̆M*d)�1m^�o䒻y��	A�qϲ�y�]��R錺�##a��Z�k��0U�%T90%����i�}cb����j��]@��?�(�B鹛}���;�{貼�?�� n��Ji���W�8����ng�;/q_����Z*�Q�@&\�������/�=/=�A��6���)|RE�Q�s�|�X���챾h|Z�K���o�h��e�+�i����g�Z����_F�]��s�-��I��y��aZ5߼o���?��	Hz8�c9Yd�8�!1�~j�� 4ُ*��	E���RI
#�LZ�!���
�u��������N��Z>���n|O���u�2�=f�RvD��!$�hl� .vx]c��U����O���H{r�6S�jh�nJ�u�g�%5ԏ�M#�ڂ���>����Y�|�m�|lt��s�6��xi8��[�w�����f�p��Ś�Z�A������+֌�Y��z�*cY
S��,��!7n�p��d� ������6�s-R$�<���A�<�o��,/���~�c�1L�tD_�B�����A=��zd��� K�'�sz���D�9=މ��G
��L�I%i����^���NT�-f-b���1�.��"@��IyN�`W�������(Iowu��D�qɭ;��jq��xG4z�-�>�C�s��ن���U�.<�E���s�_|6Ї�Ʊ�	���W��Y��l@j	���hF�b<pg6�V�[ۮP&�����~�w�!�0�1Ђ���8�Q�4�0ئ\�Mg���'_�=��>���]Y��������N��6(����$��?�]wu���P9>Nk�n#��-���0;���qɂ'9��z�-�}�`�:��lW�|�_A�<��Q���@��H�N�_G|�l?55�!qX5	�>�b%kM(��M8��T��[*��o� bsvn���4^苐 �q��)}�0,G������k��5�~9UxGt���1r��G{k�g3�H��9J���ӛ_Ћ��/gm��t`�ӯ���]������f<�	*�v����sH�"9][�ZTV�\&������J�`N�e�V��!��>�0�����a�NH]X��zF���CpSѧo�r�z#,�Bv�V8"�6��ݦ])�!c�3|���wZ�1�Z���ovg�$s��	��M�2p��,t�[%ڲ��oB� �@(G	��E���%�o�8B��b�i ��msWZZ.&���<W�k�Y.�����	6ۓ�vaB��(�<xvQ/���5� FT/�x)dג��u7���ʲ~�,�;/:�{^��u����\��Rb�)���?aX���/�8m�o���.�Ks�$�pE�</��.��i��{�tn��ۃ�Q��rp9f�Ȗ[�Y�oOo��Ҵ�]�-+�Q?{>z�]�����1G�u��;b�� �V������gV6q���&�Dye��5)U��J<{?A����߳���=�Ɇ�gU�H�8U핉I�M�P���/Y �om��M[J��ꮕD������:�~�Mڛ��@zQ�e�v��'�3�_lx�� C�,�8������qp��qH��n6�@��:��&��ԉ��q�6F���<�IX��%��MDL���������m�������e�S9Y}}�憕]3�IL�-��_"��y��,H�3�Oʇ�-�E�ˎ*�2>��1�|DANPgZx���hne�3���Nj��j����~��F�E@E���'6����fi���m"z��zI;�����65`5o�ԯx�(��{�B��?�����$��W/O�RO.�Ap�� �Å�����+(����1ˢ�k/r�٣g��FS�OO�.qؐ��!)�U��O:dE[{Hsā������w�L�Wgn|~'a��Y1k�N�D��<'A��I�����^�8˛�
�1?�!����Pf��A�K�l���Q~;��ڡ����{���af4���;�� k��Y�IBGHSXO��	�;�+2��e���Ph�B�.*z��������@$�a�����\m���{�4���Y����d>Q��~.��Md�3(p�(�$�A����}�݁l���`Ȉ��țJ36����2�������<�$�-p�ʴ�]�>��u�<Щ�Vt�Z�`��a�T�H0��.<j�`%��!Ȩ/_�����`�y���%DR��ؗ?��e��d�7-����ۣɀ����:�?����y��4�����h-����`� �,ge���"!u�7����,Hl�#�_�6�6�I_���-�ʡ_�7z5���]xBR1X�S��x&s-	���\ X
��H�"/m�mF�:��6�1�^F5�g6�4�B��	`��B��ԏ0�z�H��pO̗q��\L)�����]@h#k��"AĪ�$�_�B��G5Hmډy�ӊ��z�\�����zm슱+$�B\���3�F��5L$X�|��Y�<Ӈ�����F��G]�3�vdΪne�:!�V����sE��F�1��|*@ń�J��8�z�J����qnK��t=����_${_��{~�K��>��H�;��/���,x�}����bf��� �f�� .���?v�v=a�9n��O�)���4�쿐U7�$�^J��Z�J{��8{�I0��.��c|�S�A��L�a�|��YHא��I��~P�V���������U	zOC16��5k*���4-3�r����T�/��:�m�h���s�!����<�J��6���R�I
Bx��LM@8�D�@�	��u��t6e�k�p�ፒ�e�,w	ڤ�(����_�Q��T��7{�w�ͼ�W���@f���%�SLn
��/OM��3�G �� �Q��v�� 6U�㬥���ƶ���V�t@�X�8��Z(���*S)��ls��ݜGN��	*�AWT���W�R�6�dX.E���z�n�c�y�*~�Mt��@��?ٜ
�X�W�E���x!	͡zwuAe�]�T[�̲�kemx�� yw9$&�И���C�N�:�&��o=����e+�aH�L%�]�28WK�7��Ǡ��G��H���M������3gƿy�w}zCaOy�*,�����G�۵������sk|Ɯ�&\ňZ� �|B��+�f���qI�[��qN��;�P	D�￈�N��t��)��b!�t��;�-_�]2��&����Ğ�SS� Mr���+��nX��ء�x8�uMM�t-ĽT�����z����Α��!��8X.j�;܎�g.��J�߿�>������k%dX��4��H@��ٳ芵T�Ԩ�� �M��%���,��qvy]�r���0U'�j�4�N'��<b�}|��~z"s���7޳��A��4PŪ�nX\4�U�/
F�:C*~��:�2�r���sl�/ҷ��P2t,��j_��O�	J�I�#�N�I�������>x|W@��n�ST�da�DZur/���.c�x�����OW�ݎT����1v��P���ul���GWe�9L��tr2��M�K|�<�r �~�Q���T��[�O�a��"���J�p�x��b,m��4�M{�ǅ�6sr�[�AlT�#|J��wZ�X`Y�o���'ܯ���'������Z.� ��FU{���.m�d̮`,a���V����Q�� �`����>��X��o�L���l><G�5���
��!gS��  ��n�qϢ�����="�'��3�
�O�(e���=�;z$�|S�F� �Ǟc�E��K�G�^�!^��0���v���#�T�W{!Xk�X�'s��i�릥�g?��nͪ���x���� �+ng���+��������S����]�,ڭ���j�o��֔�o���i}�o�0;<�k�x��a@��V�կ}'?��_�;�5G��ɻ��2�ym�n;Y��1+K�|k�k�1.� �g\
e����t�p���^!����؃�6�n��o�k�	x����q�MJ�J�h#s�,Y�=�WҴ ����C���͚2
�d�g���L;���x3J��<���~RQ׳���-�.]?l.'��l��z�̋b����ǉ��ǡ崓 ;L:Z�"B`��H^Ibbw��#+�ii'$OW��~�P�%����WD�� ��ʛ��.��14�)�ĄW�s�"�wJ�6(��ρd�Q�QKI7��c�CD�J46�֦�G�$'���S��;FO揳�$�`��Î�ZQ�&��߆2.�j�ua�ڃ�P,������9)�LV7]ZY���.�G����!�h/��J0.�i�c�9A<���5�����C�#Q&����d �ٕ����Ǩ�6�L�QuK4֦DP��%�}���J#�?d�D�1�gP}��	���$�[:���0z�2��}w�t����7π���qn��%,�?�a��4n�Z�mۇ4>�^F�'rܷQ�('�8��d�F%�͗��?N9[�If@�7yyy��Wَ�w��$��f ��! <S�!������I�ҿl*�]��������e���N�ܞ��˔n�֐��#&�w��ӻ�h�dk)f�"���_H��;�
2wU�}G�ۜ�V���z���[�7s[�'���7�JzY��� tz�##R���4L�������9;�@�
�Uc�'��j�4i[�J|��ow��ט\vObi�)_�9���5(#,�@���H�a��|8��}� ����?��b�a�|ԭ�j��׵)��FF�6nO�~s8x�L���<�4�a�U:����V;H��J�e��&�c��\�k�&39O4O�0I�9Ӥ9��ZQg0�Y`e�V����\���ʠy�:�F+>lC�(��hX���.[[i}�/(�ieb�P���VُSTiq$�o�B�t~[�-�H굕��#+�d�67��{Ki$e%��:X�|���U��¨$���$�l���+C�W�0詍,��C��Xb�
��U����}5ǅ�D�U~�b!����H��mn���rs�.0}���G�b���{��T���l��}c�/����r�6��ɥ����X�b��N%��'^l������x>�����a��Ī�� ���KT�_�sC$��!�a��X�"k$�R$(�Oޘ�hw=���N�v�3*��7�ggg�z�Ld���G�	;�=<>f��'ѱp1��%ݽ�2��&���6����\�s=^��k�=����*������b¬��C0��T";ayӨU����P�ry�M�g�{�����8.�X�0���Ź~� "W�ӐzIcv���"enO��F�MJ��6���'"m+�6�I�ʝBBنq���fI����W�!rHL46s�ҥ�"�N�N$UGUX0��BR�eW0�Ø����X��j�3;h�U�Y=@��!�6ɗ��vb���Ga�+�,�sh����s��oN����i��h~��C���:�<�-q<վ�RK�GR>�ï
S�/	5�' ���^�hW�c9�-�j.��)j��ߵ�9�׾2Y���i�ba�Y�����")I� j�>� �����/�b����s�b�A���ss��ͻAN���A(��J�	D�w�H <�-������[�v6$�ԳP��bb�"���Nu�P&+��7:äN��tO�����V'�Wq#2�����������7?�k0������5�j2*��l��Ώo�	���Rߌ��1�~�ʭ���J���ջ�P2=r�΄����$��k��BC�:�ߨ �fRkM߬}~#��n1����B̡U�7�Ri��E2�e�$�S�ХJԸL+�@�{�)��$���`���J�?�s��07]5*�
O{Zz��E7|�ٻGł7N�ES_zf�E1x�$#���/,�Tv����(�Z���� By�N��>���S����C� =��>���;����q'C�첰���L��z#�kY��3��Y�E_`��W%&�&I�p�������cDR03��1��W<��o���g��<1����?�-,(�������"��~s,I�QL�-��IقKG�ʛ���1U^��j�ط�N7��Au���NH�@�K�:��)o��ђ���~��U�@�ϠK#��VG�Q|�k�C��G�=x�e֡��{s�کW��p Ջ��}�7�g�;\>F�h1`�S!�Vaƹ�T��f�a���`r�ʈ;|	h�_����Ꙟ?�&FH�C+!ja[4�R�%�T�����]���&��X8	j����F谌aF�娞�hC���K�$7ֲ�F��X�t����{�e����hЉW�:+J,ٙ#�,�k8|%Q־.e�ÐK�+)!�^
_�ǳ\d� J�xH��&����a���I�
����S�B$�z3���WJ++�ۗ�&�.~�
�<w|cT�J� ��m<�ŋ��5�:�A�O91S	�H�g��v�Ox�"�݊��\��U`��l֙pL�D��^Gp�<�3r)��S���۟��#����ѓ�3l��v�!�,�k$N�ڐ����b���g.2�(�0����>�T�W��eȘ������V1�;����z��		@#���Ӂ-�cR��a�}^�����W��GS�� �>,lq$��LQ���KӽCh �ҔN	8�T�h�a:��`7{������Ʀ7;K�1�ĎH��,mBji��Ja�����RIBߦ*^ʹF4�6~/y�X,[��R�FXJ�J��&�ވ�
�`�����G+���ll��h/�ޅ(�ұ���Q&9O,YTTFv�;g��p
��:�$��y�Y� RRip�2��t!.��'8�7��;v�7ʽ"��B������!l�?c�^�szI�"��!��!.&���ۙ=�ê���ly�RR��S�;�%��xt�������@�T�Ul������@�"�)�.@�I��m%	�e�J㓕Fl��eH$^�����b�~�8f؁�dcLc��Qo<��o��V���eM��K|O�l�X�����|G���&��l�΂�D�M�h,Q�`b��̀���5�v�f2��`e����R�Y�mL�)dM���R��E��Ƞo���_T��3�l]ǖ�
C�Cm�O�QC ��2{u��F���*���� �]���4�)�l�l��u��mm�VE���\��q��${��Q]�t��������u�������Er��R����rt��ɾJh�R�����L�1E���bl�0�jsL���H*�L�,��Vsr�z֢�i���{�S�����b����!nb���E��v�.s貦�q�go�#?�t�h2b��H}� �|e%D5ȃ��T�e������^���t�'�)���������Or�D�0'���2�O$��{S�J.#~��h�ុ���񉧑���K��u��~�Ѓ�|���@��Y�Dk�Q�m���"�lH�z�|����w��T��%/�!g�EX�w��� E�V�]��jC��c�s�;&�EUk��S?^k����o:Y�<��ޡ�88�;�L��D�K�������X�oc��P�B��Vzms�֒O$v�$�Oys8�\��l� �������A���x�A.R4�s������E7q���� �R��w���ޠe !g@��6�X�������̥�*��>\;�������m<��ޏP�=���0���9|�A�ڴ�)�L��qя�z�^,+�[t�|����"��E���[&��^���#�� ���6r����s�o+�޲|��>�9�m�_�tv̈2�ۿ�~��K���3M�D;Bx�8�!D���h2Qf�O[�O�������+MF���3�O�S={�=3���P��['�����L���ug����M�����Ue5[�P|v_��A3�7e����)�w�` �xT'K�ID�ܐQ�I%R����A37�%|b���DU�i2|�Bf��]���BW�<-w���ImWEd��?�@�r	:�r̔�!�k��~�;���Q4#���\dG����d+����y����J�,C��"qL$�f���cB��`W��m0>S�8���3Y��d�q�O�ӌ]�z�`g&$,�rbA^��[�']�Lr͇k����O��O�Z��V�ꏙ��X��?������Z.ę��iS�hV���3�T��81���V����+�h�m�[vO}����<��otC&w�-a�2�K겢`d6M�� ��g�B+K�>�հ��8E
�ln�XR	��`�M���|R�P)�+|�#M�k�țT��0���iN������c�P6�$%-]�G��QUZ���yl6T�&$m��TȮ�K�L]�d{��`U�����q�!F����{��R��x��5P������ڰ�I=����@^V4]������RnD�n-j�7��%�DQ"_�&�҃5p@�r���Ԍdn�����cW����d��O��W�K�`��Mi���N�����K���O�K��_��&�I>�R��A����q����[����F_3c�G�V\���#��Y���*9�F`�m0�q+�Z|'��9ЅQ�(¿�h���[э��%�ȴ�j@/��E�����L�ݦ|r��}���&A&��!T�ecF�fG|~��M���.�>�%�����m��hfTusn�%�o�W����,���79	F�%N�\�ϕͭ��
�(�<��~�;,Z�%r�I.����2�9sу8�(�W&��s.��س����+�1��Z���X^��מF����X;�Cq������~Z�!��^�kB?����q񀂕f����k�G�Rfܴ��o�.�鬒Z���V�"�J�Ҭ���i���Ft�7�U�R���5d+����@�]C̞0�a�Ѡi��lw4��4J0�O7�����ntw�����Щ;��}3��(�o���P-{1c�u�du{�=Z�<�ظY+>D�W��mϖ)�I�*�~�1��	��������8��.J�UCPkk�˺>w�4���KQ�wڑ�n���^��U�Ym���~�b�����kvGV�����E��z��
-�
�|\��Č�	g��c���%�Zk/lR��s��KZY��w��mƏ��<��*Ϭ��KD ���ѹ�R��`>\V}B��1C����a�y�J���ң�&\w�b��8<)�ܥTJֺ0Yg'N��]F�S?Z�}�%�c��,"M�2�Ԃ�uM��ߊ=X.y���T�����V93٭�h����i�7���W�X��^�	Bi�J�cK	�>WqU�����n�9s�.tU�\q�P#"	��Ҹ�,[�vg0�x�����,��g|xDV��V�ť�Ĥ�}�ⶂ�ƅ`��'�Ɛ�xu�uHG��1��#;��\��eH$���˔&�҄M-��7�L4c<��9�h�E�@���ʭ�ꐜd���[�z��h�9j��;�L��;�?�H���`ȆlJ��d#��j�&���}�M4t�����K�J<48N�XT��TZEB��~6�(yo��$�Izg���I��g^Q����I
0%�fn���CL��IM�z�{��%�^fBA���ư,��[���ُ1�P�o����9�
�ȕr�q��3��zF5����;��cޫEfp��MH��nK����ޚ��:^]�O2��#*�����-�$W�lO�l�Z]���F���a-�rxJ��E�/j;��3ʉ^�f;�a#:�iAuЎ4�4\�Y_8^�mă�Ӗ��n�,^��΢�}����*��ٮ��*�`�YwVP�X�R(�mڪ8���s=#��!.��d�y�7�:�����h�s e�7h�oLL��<T���v��,:Lf�kM�M�o�I&q=���	�,[=x��/�r/��9q��	X8F�o���]}��_�yDC�~���5y:��\O�{�u"7�j�0�� K�52�,R&��*�����.��#�ˍN�K	�=u�?�AG��M�j�pZZT(r�>��n�.|mYJ(�b���E|��z*�,[�v��-�-+��on�*%|ߊ��#��6 �� ����%(�NJ�>�.[o�R�/d嫴���Er�j݀Ҿj����F[�r�I�uG���׮�7�@���Q�V�!��L:�C^���� �i"����אF����8m�� ����ShAm�5������O��<�����?��I���T��Ȫ����!��E)�Y�9J
�����M��X_��|�&�ȸg��O�K@��#W=���x������+�nY6M�徟9Z�X��X�B֭зg�����`�.f�k2M\Ϩ��F�Js���#�X�8߃̯,�[iN�=�h�C��9��5��1]Z�B�m�=L��ޝuՄ爁=�:�'|�'.�4����Fo��v{41���IW�YO���\��{�I��������DvON�X���"��(@eC-�8UW>k��:�&�ZXZ��L1jYn�A!�G�<̮�A��Dj�%�@��yڒ�	���P��_����0.ɘ�k�U���c�_r��� :��MZ���L�#�B�r:�.���̔�ow-���rw�Z�r�ȹ�u��}��m�\{r���I��)7.z\\�#��Xr��2^��3|T���7���d.ԋ�s��cI������Xض��qv-�}�too�Է�Zv��������5~ܘ?W��Ċ�#�ˢ�ĦX��ޟy�����=OS�����1�K�*ʱUQ���+RzY�����'��l6�ISN�ј��ŧ�)�����{ַ�;vο�-��y֏'v����g��h]�� ie6I����������ǡ�1�O���;w0Wl�0P8��Ӽb�]�e�ήv,�5I��>�׾`��S�l����9q������A��y�Wu���v?���k�������vm(:�����i�	q_*|2f��wg����7���M�z�������rI%iY������k}U�k~c��ٽj�y�ީE��v닷�n~��ǥ��^�qt�D�ˡ��m�_�~�������z��\��������lE��
���-����i�=�G+�+���w�<͠V��oye���Ck��Ņ^���_.�{���/��#U�b��j;��s�����RZ�.:�my��Hg�����^�䏻.�m�l�_|_��S������|�������oI����7=�n�u����_,��P�ܟ%)��!���h��N�,`ë۟k��T`l�U�N�3���jȂ�S�⼁�3�L׃�3�κD3��f��v��l+�I1�sԨ��W����n� �־�(�Am�N}��C�f}`b�B�;�v	Ƌ�ME�����:��& PK   �rZ�^X�� j( /   images/cfd750a9-6fd4-4ac0-902f-08baa65eb73b.png�wT���.u�Q0@�hpl �Ho�p AA�K�#�?j�q��RD� ]@�Q)��������9q�3�����{ג�fe�y�����~�y�p혁���«	��_����g?��U���z����y��?�OЏgi��O�G�=	��e�Ο0�77{i�y����=}�����+}�������������j��V¯�_N�Ų?f��[�`\]g5�Ʌ����+�O��
�J�[��	��e����bC_�6a���B��OFu�;�����-�K����O�|����5���m�P۲��vD�ي���;ŝ翿m}�?6�����7�����o�}��~�����7�����o�}��~�����7�?��������s�!	�ʁ>y������	�7�q��bu����ecɔ�V��߸������{d�g���W�<��B���I��[w�u�e���rO�w����U�?}T_�ʰs��%^K��y���z�0뎈�7[�-��=����Ȼ��;¿�O$~�w~��������< �������� |�����7�oӔq������|9�x�oד�2Ӏѽ�Zd�6N��L��ܥ�X�r�?�(�geV�n��T�
B���+�ϝ��w�_��-���A �O���_ �o�}���6u����p~��V��-J̞�Kah���L?�Y�/Z����6�۷)-��LMm 7��5�A�q�=_U94bj���J00d.S�*�T��T�ɜaڼ����6T��ŤÁ­ڝ�JԥyVAu�S?�K�H��",ݢ�zx�d�&�f������I^��G&t�+�gE�p��/	Ji�$�N��R-�n��m��!�������X�T��dt &���;�Qq���xx�.�h�
�������`	�|���fG�af:��-��1�C�Jg�/VO9�f�WwY��|�:���I?)	�Jg�(��l06=3��.V����z[��lM0*��[�㩕c�SmnZ�eoz��[��JUիO�:�|o3������(V\�:�g�㠇��kU�*׀{�~�ME�Ϸ|@0샵OF�X����Mi�S��N�J�HU�j��7�do]���5;6�� X$���⯷<;�w�t�b���ۗ�9�iȀ��g��v$c=�7sՍ�ml4��?�ȦUvvɉ��l~�|���7��VUiFA�Q���]�i�*�.�8�๺���-O�@ol���a��Kg��5���R�p��I��4N�:�x����/kV]Jg�f$5Z]dbbi�����)�٪A��3����s�bu+���41�5)�W(���!EEE?u��M%��n!��5��߮隗d��+�h�uF�z�_#8X�<�@�[+=eҸr�|[[�-?�%�O��I��M>����>�̦��<=�/�:׹���o�����a+�*���\V%�����i�[�ZP ]���KE��Xå�F�5��	��?�b !{���Z��Բ�����������/,�����/�m�0�'������Jvkf�
��楐Q���j���J�����s�3KA;�������rc,r� yC��ξ�����g����Y ����(<*D��P���4�U,M^�hؼ��������|	���Z`�?��[��k{cen�
݉_E(�C^�;l���,.���B!��r����-Q����+#=���8mE���3u8 <��u8;^tb�õ ��u���b�$�'v�
��� �C�M���<lt�b_z�u�PZ}-��'w!����bA��n-���̌�ig�P�(�.�o<�`2y*���n����F���H��	*K�ոp�������~f{G���%��7uWΑ���'����,Rw��ȐO�θFxFU�tb,��v�.,~���&4�Y����Pyee��'�8'���8�=�%gsW�)�+\���IgU6� ��o���d��_�c�o����X٣�r���My�j���9ڿ���.���S���,@�p0�J* �0*A���&�@��9񲉹���t�e�'a��b%L&���-��`%7�ǐ�#SҹS%�r���X·��~��h~{�M���������l�P:۹�)��K���H�D$M���K��HI��|y�E�K=��\��i�0�����~�|�9B����ۂ�j������OSSP.  �05��
��#���3ǥ`�w� �-[����>z�������Y=��Zf%J�\bxFJ�s�?���C�L~�M��b��G"�RS�CYN�=zqTҸ��ǅZ���7�!T���pj�`�����woI����BB�/�*��ܴ��	��XO�I���p�sZ�o�H	o2Eh���?Ǽj7=-��#0�|�%G����}��$��.-�Y�Z����I��s!�K���=:drQ{8 �9���-7���r���
ée� K�����k����:�$���D����Ԙ��_�W���T��L�R`��� �ek+��� �o�&猇Ǿ>����'(��;��/(Y�|W�޷<�a��S2b��lM��]��X��3�o�e�;t��m|���P��ܩ9�l{��)//o�=3\��B��▣�c��Ϸ+�Q��@��r�FMxͪ���?�P�a��`�C�n.�޼�}s�/ �;۰�'pc}�l0�hqv~~~�2��t����F�u�^g����S�؈����9���ts��{�5�gS�\�B�Sf�Fv� �yZ���Y�����>8��|,`#�� ��������G����	����� av��2+�~Ǡ�;8��e�P�-��-��[����+҃�&K �ʬ���&ryP�5,�=�@����d�DEOUDH��Vd�\�z��*�h���FذC��Aca��Ht{���;P)�ϟt���t����5Q��n��K&�,�k���As��f}�^�Uob7<�Tc�:"�)\C[E���u���0��dk���I���Z�rS#�d�`���b��K�{d����WW��dI��%M�n�3߆����w��V����P����'����tW��fL%ߙd�ژl�'����N�7/���1A�,���
�"w����n��Wh~��bR/�oڣT���+�F9��Pǵ0Cs�l$�^ x�-}pv�6I�;��������x@X��4��Ѡ���8��"�ͺ��1��I݉wޯ�M�z��I1u�S(��׼G�^\.	�*-�\ �}�Mo�+¿l��A["�7p1r�mQ�1�t"�J�d���ѽ,���H��8��TI�XCg��Ź�N)�[�̙�ڪ�]�:K�3�,
t�] �W��n��b�3RN�5�Ώ�T�Y��3��*((������w�:�n�i�M(c�{�Hb)/�666.��s�ȝ"JH�Ȕm��W�\�}���(�K]G��߭~�i�RZZK�in�@��ѽ��\�����[Ce���u��⩎���Ea��>�r�E���O�t�df�\��n�(�_���!u78����n��H���Mo%u%f��@���t�&�k�ĩ��.j��ja�s�T���?I5%u��x���@
j�4Y-�s�eww���6Of׭�ܱ�ySuu���nQ��Bm�� ��U�5���1�"A�:?=���ّ��y��ݵ@ų�m:x�v���'��뛵ʛ�tw�&X��τq�z��Wҭ�$t�$�彭;�T~�\t��xw��O�g�=22���D�C}��z��䠑.�;�8���>�Yg8�X�urįU��� ��q�h[�^�4��*�C���s�81}
�AC^���f|� �j����$R*A��L�$Y\�	�ɶ$2S>Ul����k��w,�\�ׯ_�*�
��#��G�����ı��;�}P4[v �C7�>}�4�ݵ̼���auab2|ƭt��j!����5KDɄQ ^d�^em1le��!�����l��-~��%�ׂN {r�0���Z5ab�M��H���6�в�̌�����90��H�m���j��vS<E��Y\CpmR��ݻW� ���s�&q�)�� ��6})5U�yN��^�_t�𾍴��^\��Qq�!��^�<E��p�b���{G��q(�,3�[�ѹ��A+��`�0�Is�P����=Q��au_�q��I�����zC��r^�Bw�y���������d����r���?��Lkg�یp*���m�hL�U�n���wq�}�HK~8�� ��.�N�||G�yv��ݹᢑk唓8^]*8�<�^�z֎\�Y�b�����=��_S˖.OLL��+WV/h�$��vh�U�ye�H}��	����Xͼ��Yw�g�>����5ޕ�w=��}3�����6G�v���ќ�s�����E���D{��8kT�M�#v�f���+f�V\�8 �o��b���៩���c���%uGP83��t�'
j��S�?1fb�pC|�;<8%--]����8����*}���H�fō>��P�wC>ir��m��
�HTy��T�O�@cG���
O�XZ���#Z����}s���l�'w?��V��6m�!Q�����9������qOM��?�u�uC;	zL����$�~ҦΒcSS���z���0Յ��z���� ��{ٓ�UI���]1*!Db�m��!�/n\\�j>���-3�"]�Bm� Q�Tv��n�|�8{ M�N���ؗ�O��Y>*qp	�D� 7��>j���Y��`�4+?��F�#@s�x}111٫U^$�}�} jõ�ڴ�I��G�*1&0�Rv�hM_61Y�M���q��Pv�<�1MM����1���#TIh����)ɵg��g�i~��X��#�n�n{['�AJpJ�ӱl�Q����(����4ItWЧ�Y��w�K�O5M$���2#��Ex`�P��zyS��/кI��ť���j�9��jY4U�����'e�	}~��,�pp���\������q��(鄋�X7�������%x��e�8v�f���]n��w���5�/�MML�6˄���X�s�N��iD�'�A]�\�԰��U�k�"�Ϯ߯��8�I��7o�_ᅅ��A	��T2{/6�"�9��Ѭ���T��'���q�n����K\����g�9l��Y�$k��j�*��6TV��Yǭ��c��C��������#�.Ǉ��	a����k���P��H�*,N��)�C�XF$2e���a��D�A''�L*6�%�5 D�-���G��?i �+�;�Fc�J<�fcQv�4MX�}k�b7h��c��D��	@y4x/�}r���	�R'��h�]��L@�n���:7Yi���)���6�,5�ㅷ�q�ad�؁��4�-F3�ƅ!oʊ-[O��� �
�P�^(Ij�1�6Y�����X�������J�ĭ���W�ֲ�qh��]Z5@Y�^������C�_�&Q�3���2�q�>�^�- g�[����b�
��E���7������m|�Ĉ�(&�����5I\��\xtgq����b	t��dl��
-���w�ܮъ�u3y�V2�'u������w�ݨ�}�,,\��A"#ϟ�bX�~�X�jj�ujƵ@U
���T��b5q���,7¹W6��P%Y� P�x}�D�\�_����f����̑���%,zD_%:�Tb�mO*�h3�מ��W��=s�CsA��\�M��2f�U~�E�ͮ��) 5��A���F*�8;O"��~3g�2�<�[����)7	���~�Nׂ�
�i�CEW�ɉ���j�c��J|ROW!-n%-� �q=h���x#e��̲a*/���<�ƒ�H�ґ�ڲ���e�?[�q�H���[U�����E��[jkw����c�a+E'e�,;nk�mU����_�\3�r�؟5�l�rV���+�������
��/�����먳��O��{;���ӯLͱ��S�fG�Sy�����||'����� ���utt�\}��/y�L6���T8M0&(c]�鍜t�C5ɐnjm�K��2P�;P��B��1a4�;�t����,�G�H��mF�a�t���ׯ_���aߥM���E��L�u�h�7nܘ7����엕u��"}ь��\~����Ke�ř����U<<i)���<�>�J�J��l�R�_��d�݃�.�\��x�yP�}���(��9�����)5Pru��v��h�>ٯ����T���'[��{��B5�z�Ʀ�����m�Xܧ�[�ǝ�i~�'�,t{2�}%p�2�m�����رsg�\uLf2��1��]�I�ZQve�jj����m���֮Y����<��9�L�߿a^����_�n�o��$�X���W��D5&0��1v�0������2�ċOJ��.Z�$9��m�B�*����!ذ�� 1��kp�V4��>w���}}=�����%�/��$O_y�Q�`r>�
J�顀f��$;�^�xq)�"]C��)N��M�%�&���@��]f�5i?6��}SӔ(d�,y>�a/�t�4&�i�͛�w�h2N�EԖu�}�v�]��v&G���%OZ4ɳ-v��r��0׬��������=�#	V�!�\Lwe�%��d���D�m`6��,B��U���į�<�=�x4�� ,*�`4?����P�=�?v,��?���g��hI�.����_lIII�)
����P�^���k�����@X�x���۾���4M?ik�3���(�'�ӢT�x|�ƇfR�!�V�:Q%�z�f�� J2�A�.��S����!΀%�@�O!����фh�Y�"��5]�z���)'Z�W�����G�Ç$:kMmt��_��?dT�?ލ�xP�d���'��R����{���h�3��f����R6��Q.T1�qc�ܙ�Q_�Ŗ3�Bg��ҍΚ���g���D�,��b�oJUkee���L�<i�Z����Af�9�n$�&~��EQ,��͛5c3���ib�")e�^؍�0hnn����g��_��y]ݻ+R�~��洙�@��tH{BمP~BV�>�<"y�H��SQ���p��@���ԋ]A=�����~�+_@��_1aJ���ۓ���)Z�)�Rӯ�������_#P��q>P���[�����v��ʖ�7h��L�L������`�͜���O6��rˮ%�r�_{4s�"u�ԔuA��U�oo�`�'Rc�93�U���4��:"��ȓ�i�����	�^�fvNNΌe�`z��ӆ�6�>ni�$,,�{����	Y���)j��Cۼ��4�j�_v̛M������>+sb|<�3�l� 9Ȇ��JQӥ�ُ-�dd���ɓ'����,N�.��Ӝ�:���:ooo�_������uD���������0��`�νg0&i��Z�WY����L������_֣��Ba�٥��3��g�x�#�����:�Ť��E��<|�V���Èc3 /y5� U��s��$�y��8��6}?Œ:P�4Ĭ�Bzm���E��#���9���.I����4��\A ������ D�3(lޒ����c��v�O�� ��Ņ�yI<!����T6tn��33�S����ɍ�Е�7
Q}�U�8P#`��"���QBs=�Ni�E:u�TU�gy�z���
3+����f�����Ͽ���0�DW׽{��?SRZJ��VR��?&c�hӇ��4�4F��m��o���JkZ�Q�RO��?<a���bf֊я��W�&&nV���;�'�h�rB��<��<���狫�Y^�Űdd)
Z��+C��� Jv궹KL��w.g��ￚ�陂y��x��!KRJ���Q[����?̉�ݍ��������ɞ�?��GP�}�F�mM�_�������>tw�(�Q�.�����C�ѝ�!<��N�H6P+cm�̣Xl���Ѐ����g8!{H���RM��k�����o�li������%�~��6~��줱z�a5a�þ�(�|���|OV�˧����!�����'S8�{|����Z.fE��ф٣�q
������ E.?�g��p�Wps���<Fj|�R��?��!4 �GEG�R�}}}
��RRd�ѯq<i�]�Wx�v�P��r���I������\\\��ik`"�~���	�� �	E�f��},��L��PvQ%��$p�r�����W�*_}��!�-L`o�ʑ�� :h����q+�K�<�M�aԊ��O.u�9���� ������Օ#<7?$���>3p��w�nt�st�B��ĭ"5z��?~�7c�죌+up��#����9�nu��V>���ciq!�����gYY�"uK�S�R���.D��Z����C�b��(���9��w��9b�3�p���N�|�!�_�=�~�U���f�8�~F��эv�	=z�
Aт��oNɰ7��?L�� ��+p��GAff����� �d�A��&p��H�q?B�i�Z��8.��k][[1D���k�WYK�	�b��ե�d��?����啔����N����S��e��_�8�n�6��'��&��.ED�O����!������1x���\������@�?�2��zP�t���acR7�ԣJ���/��J�����(	�F$��@3�	c[���?��ގ���?K;�a~��č4����r: `6��3�C;
��Rt"��Y��mmm%����1mYF�ݽq5:VAF��G/)'t�{���4�����	�{~ε	�K�Rs~����|�׵�������3�Oo�j������	���� 
�%��ڐ�){���a�G?%&&j�F��ǉ�Z�\>�ɘ8&h\ +��2%�=1�U�l�~n��!v�&-$ʮŐBz/��]�p0P8w��6�'Vͪ��WE��1�Q�}4n%�Mv̧�<�2�7"��J����n�	�<F�0��bJ5蜸�rد�c����A$�i��o񰰰�\#�LL<�����Q�����2�+3�VoooB�˂}ƈ��p_��`v
G"hS�d�n��5��U�g(77�
}8����:뀢�����ӧOɐ���/7�'����*�X}��v�ڙH{$�1Uv��^x�����������TU����퓓� �dgg�R�%ty�jppt��s���b�����
�jvps[�|�◥)%��QX6D<)**��>}��/�5sлn��v2pj�d �B<Zw/���4?������k�Q�xW��|҆ԝ��իhH3șh��]9���#'�4��Zn�X�\�U-J���=����s�&5D�� ��/�w[�����2�]�7��-����1��/]�k֬�oTc�1I3�pe�B�QJ��[��p������e{����|'���IӎeG~���XH	h��s�!?#��
�p{�M7���/g,"�|.��]�x���s�ǴC|MG�ǏKK5�s�d�����_*�wbD�&� \	�V�N����Mf�1{�������t������,V����@�.zA��ߺ.ԥ@��
	M��y��`�#�y^2S233���*�ar���!clu���ÓE�#@O�,?������^<�������KU��.rPl:;w�����{�%F�-��b]4�AA���f@ʈ٩S�0m���/�u��G�a��s��~����V��k��E34�+:ga!��F�	O�X�Q!k.�ɓ�o������!t��.���d{{��yyZ༈RWtɲ,y��t�E`�N�vĴk0Ӣ�@3�M��5���Bt�� ~��>���L�gF�i�嚭��'k�����B�� b�Iݶı�f���191		w��}8�,���0a�yB���͌�P��q?0�������� �p��e���������[IT5�#(�,踩��Hx�/s@bh]�]�|	�Ҧ��M���_�Ƹ�}NI�Ourp�s#�m "�on�,�ا���FN���Yz�

;>�bCc#D��뷛����אG|൘8"�� �J%a��*߀bw�_��n���T#�8�O]K�fQQQ0� 8Sn��.d5uXS5�0�ߏ{j�UH�RB�ɴ��v�(��0����~�i�l�3@*�����$H((�f����d�Q0S}���I�WB�S��Yf0#A�o�F3d	�j7Xy��dKK2p��z�䰎�����6D����e�O7�Ǉyyym��=Q��0R���J�F����#�K"�&��T^~̎��	�WaB|����9�����Sh�i)h��Ko�%��e�e�ٹ�2U&X#<P���W������?�m+	TL5YN�*@��v��f(��˷�w�ݸZs߁�8��xd�pXKV� R��7/!�	D����s��&VO�mcC�FSu�����ӏ��o�^�#Ȅ*l�Uh�����Ʀ�T5U�D�:ğ%�4��ȩU`$H	0�*�d&�mii	�ߒ�A��!�~�H�g �@�0@���o5���ΒY��
k��'���hik(�m*��III0T=<��5S��}-c�q5~5�R�RV`irsc��+��R!��,�=��(��UU=�q��ʜ�Sr(q����i\\\7eCS<`U9�m7:��^�g�ۋ�y��E+1�� \#9xEB=��lX�cz��6�ƅ�xI]��C�`y��Fo"���k���|b&Z���?��IFFey9�U�B���8.4��!`�/ס���Kzi~��""�å�u*���>bR,*��H|���u�߿?lllLH\<^�m@L�1K�- l+,���O��rQ�|�y�6ڍV<��3kh�`�(;(���P�
A5�@��u������E3�����
������%�h�xLHHXx�����>*+[����	1�Ah ĩ��9s�i���WT�k����U~�p�$��/g�i�M�S��~�Qi�VT�����~7h��Q��e>���ӃU����	�Fh���'Q:r[���uuc쮮.��T�[_�x������ ��i_@�1���8��@59Ԋ�9��ȓc��*�R
SQ-�� b�A�wA��.j��߷��i�fc��[�ˍ���������q/4������DU6ꄋ\{u�_��:Nɀ�:����Y���VBr�i�N��7��!����54� �n-p�z���jtjz�M	���$T^�/��K�#i�o��w�XB����U��~aQQ5�y0 K�4�*���A-��͛��fO�<y�00s&[��c~zL���# � ���� �����(eH��V= d~���H�c�\���N�%
��ս׃s��r�"M҉��JB��zB�HX��"�j5���'������_Ӧ_ V�������GD��?O��,�:�Zk�pik:`��S��+��їAi���x��F;9:΂�0#�)���YX\G1EUkh��gq4Z�h!J+J�ᔋ��'�3�`�0�dT�B�T���8h��E�mB����~�b=208���&�
 ���]G���mTI�*mm�E'��^�W� �Gߺ�Y�<e@ t�7T�����C�����F�dD���l۪�%%�8���$i���˂�b��u�E�b�����{�15�<�K؊Эڋ|m���\�7�������.</�u���ȠO<�y#<����ɨ���tyC�&��}�өt�.������@X��8 $�F=U�\9Lx��S~f*��ї�t��R�e��w�����՚D��5��فq�Uq_c���P@�6?���@ӎ�S:��9�B���	l�����1��B��,�$Q�cA����b�"F�ۃ����]k��!d�&~ʖ��b@��ҟy�����a�O�����z��%��kޗn�k�"����ZȖ�=P�ť�Gx`��'{�7;����H�R��C��	��e���Y6�>\vf]�ϞL}��I)dq^Q��2mZ�`�?�U��Ot?�jJZZ"i�����|�S>���IK�a�q�&�p�~��LI�9�$������qu�������n�����
z�F1&�pqM�d�����ʄ�:�(�K�dC_jDJ-�MM��/��sR���zd�o�G�-[�P5��@��;~C�a(d�_߮{�v���aO����M����a�n�0J�5S��O)���Z�ѣ�o0;���Ga���\'B�憝dtP�=���zb�I�Կ��lKt,���O'mNWPP8��������1)A�T�C`P�x�͈�q'��<�c�����#�Ǉ�Y2SSKS��64�ۯ��-��111���n�@���ΘB�&�`�Gv������a�f�
		�&��,���=	������h_"h� 5������g���Q�T���Q��2�U"��)��\:m��5{i�R�K���+�����T;s��ĝЗ�;<===f'�y�D,_��@T��r������K���S�ՉK���V�zfQ�ܑ�VTR��7/��S��������r�h;sa+����k�q�2�B$M��3�ȋ�[I��h����{��q��B�2,ұj~�!��Y*�n�@)�{�Q��z�����]۬�9ž`�.�Kk�$z��WX��(�����$���Bg/=�7�������L�q�Ô��P2�_�����e^M?�����ذ�+�,�cOz�Û�a����^ѵ�6ؔY��N�,��^�,����Њ���Z(��s����7�<y��b.UЦ�S_@�q��H~T�܂��7�C3oۙ#)���N�5ǥ`�b;���!�7����"Cq�d4�����ɡ���;��p[��
%:�E�)>��R�<�%z5�#&�1D������T�X�#��p^s��H*(��9J6*F$Q(C���?ĩl���@򋇢�3/9V��"	�Am�ڇ_�^4� P��u�<a�ʝ�2Ш���Y��m�"���k|e��W焙G��q��qbQ�EG?tv.%AQf�	�	~�sB"i��oF+�wD஍U� M���T�0��	CR�t���
��:	��*ʮL��ۛ����� ���	Ƕ�Mo������]J�G755�I[�S���X��-������3����]?���LE��������G�� �<�
琢��+g����f�`J,�A+��O;::� O	4M ǭ0�G�\X��)�=	�Ȁ�Gd�A,��NC|D+�9Gjn�1�J��H�^�Qr|@jFv��%�����'���@�7�J�I)���>�P'00m�7���wG�C���0�C�F�}�̯���B�Fă���b�@�*�{4�RU�2{�[ͣ��=ԑ�"�b�@�V�~��zN���<])'�`R�I0����̾pQU��Xt�	+EJ��i``@���[���֗(ϢA�� B�I�'����T��S%�M�6��?P$L�_�ᯄ,[{�L���(3�Z}:�%G@��cvL|i�0e�Uq%��b�`/�� �}��w�J~�a8E E: D��E��a	�z�����\�2"��:V3d1�&��X	���M���Qx��UbVޚ�}�w�{�Ɉ��pZ2�Z��Ԛ܉,+2�r1��g��y����\{�6���U��Ĳ/���v�^6j619I�O<�l#Q��9����Vg�⍛I555���J�d4	��Bjr�)h:
�XDG�O��YM��b===C�PWTc�# ��G ��D��3���^���5�9���!t?BQ�ۈ,��7�Y9�A�I��KG\CQ__��ﰕ�&U-��(�#Ү%�M�B�v��E6�l���܏���@z���Hє=3�faa!��Z!������D���dT�RRR�=|@���ZXX�μM�H^8�6m�X�p���Sԙ^�{"��Q���J�6ӏ[��h��C��GI��\x&�Pc�::�ɰz��9+�	L�0m�=���$ ��=�ОD�v�^�<�f=��Q٣Mͬ��qQ���G��X�@�2K�������ja�����2z�,��)�7��{��l�iH1��{{wWt5ؔ�&d���#�0�G 9�\�j�o;��fn���f���܁���&2&>ހk�a��n$T`d�JI�� �����[z����@�2����Е��&����,P+j��wP��~���2B�F �����Õ��VǼY_�gܓg�4JK�yC��և����eHׯy�>���(fH�mٲ�p����� *F��h�L��'%���Mll>���N�]!9s\݈�Y��):�����<��Dt��EP��#u��M���n��Y��'�H�I�㷁�j,ll"���%Ϡ)�XBr�j���B�i
�yTIhg#T�>
��O51մƁL����s�(.ϩ�{�1���OE��+*V=�du7gۢCC��)ؗtl��_���]�>v8�	P�G-D�4 ��x3�R�]$�N�5b�ZSa�Eԋ��飽�r**�L$p�8�e����'�UtwF������򚣶cǎ�j���P�뫭�H�їm��ףY�M�js��S]+	��(v��Ǡ�w'��,9����$@W���.�����q�'���Z��it�Б�boF8�����8v(�.DT�s��i����i������ ��0�Q+�����g�B��E��s��,&�0�'�	&G��� i�SU�b�auͲ�U�+ Ӳ$A˔o0T#���Ɏ����e[�/2.�
ReИ�Q�=����g�Ɔ������O�κ$^y9�x���>9����6����f�r�M�*��ł`k��}�G��2<� ����<}�]N&{"Q�M��ܤ�\v��J�ư
���f>�ߺ�B�^�*���#PG��~��JJf0��ǲi�������fz�{z�m��z.lO�ӳ[`k�ü<y0s������h��F�ao�pڃb<Cҁp�ZXYݐ4�(\��}�v=��5��n���R����)U���1[��p���q�	����#or�����ͩ�/-.L��	���������Q=��<�M�I8UM&�=���@���+V�4EKt��&�;��T@?]H\�0����?a�@�hɵOz�xx��F�ińR���F�H*�*��XcS�TS����� h�x����_?=����F ��`ʉ�h�ۆ�ƴ���/����D}�����}��	Y���D�+֧�Lۧ� `��?A�]�?�خrԋ]�-(( Z�OHUk�ut,ցv�����_l ��{Y�� ��,Х�oʰ���+�K��sЁqA��P����nW$U��)�
O �%��7tϤ�6kFBQ�,�ͯ��C��w�Z���u�������6����;`���*�p. ��]>���͆��EyMMq��7��}5�����BK����x��-����a7���sN[GG#���0\Y�]��'��E�eg&G�k�O@�(�HH�&�1w��	z53��ޮ�a:` %y :��&�O�*[/��
���ѡ�|PB�5f�"����D(!�����""�N:`�f�] �P����M�#����6Ȕ�݈�H6�_V�����MfR��ɂ%��ߵ������}t�.+l|b�D�:��x<�pe�͚Vt��T$����`M	!�Dۼy��t?&��AQQQ��t�i1ٱ_CCL�t�V��?|q������?SR~�[�6�'�����Q��͟ �K��,�4���t�5&F֙۠"u�J�'����ѭL�(Y��ɴ��O///݁�(�	�tx-_���d�X֌	M�s_�"��S�L����'�'7'�i�X~� t�3V���4��4�V�k"u�+�@����7V!h������K�s�������5����z}�S�9C�U���i���.�ۚ��ā�B�xzf�cr�`���T�6L�<s�d�NW�ʐ:k�O��_P�'�@�f��F�h�~cZ�^RR���V�zřX����D��R�c��_����*��/��-���s@�2�z2M_ȩ�8��ـ;���ɂ-�+"�F�-�-U�	V��"�}�R�&���%������UfY����m?,_�|M�ژ�
AV���G�n�������-�k��0�ynG\�zѽ\9�s��m���������w����h��q}}��_R�׬���o+�������ş{�/�����#|i�#^�4�Yy��Țք��!11��$(������-y�<�����l�U�	�$|(@YL::�'�'�.�$LP�x����4�E�ԟj�4|bS�108�M�F��X:��4� ��������^u>�&Ұa��j�����Dnw��V��p7�Igq����^G]
��4x��2ce�Ȱ��@����1�mFf�����Ö #�s����_�M�z(��?�uF�?ڡ�����1�a\z+r�����fj,�uJ��H��/|��1����@�6(���A���4�˿B]�=�M a�>�n���Ók���Wǰ�|(�������SAAU���]}=�P��F�l2 F9�-�Б��D�Ra��7���Z{�If�Ǐ脄�����_oEHm_���_�CۏƝ�C���� �]$gL�NV��]�~Q���n�/^���+�G%�� Ł�UP��x���'�W�/^l��Hv��{�2���n�����g�8���0��Z$(�\�t�x$�c1úH��>e5>9�sm����铙�D�N�������T55/=}�/�-�SL�� ����n�� ���������
��@TAtzJ���:��������b�W�nD&n�0Z�M�8�?A�������a�HrF�h����@h1?��L?��"����!P�l�s����lj9�K�h���JJB�l�WP����J�|nnQ�l��SY�|%W���Ç��ȹ�rȹV��ŲL��|�62�����hr�G�����Z��o����&@7Xv.�o�]A����� 1%�<L{ f7��RN�	�m�PP���H�2K���B�v6��YE�C��;��^��w��=kBG�kd�Bp{�����3	K���ϴ��e����Y���=??��)UC�#����;o�B~��Q�$<Y��$�On=�>k. y�	mb��
�{���������ɰzt��q��Օ����v���q���=]��
��p�uB�og�� K�{�}[�(Q(��s�Ǯ�1�OQ�����(PgDb�V���j�Xv�qp`#�ލ74���PśHI���.{�i
�y�4x���=����B���b. ������$�4MGG�`?�S�yb]���ՅemQj��(]z���������p>�@����3�
���� �lv��,fW�~Y�vm6ua�:��Fʽ79�H���ւ�Bh
��N��yW����q��7�����pmSSS4����m��?�̲�*�|�&�W7n��a�|YHgi��Jb$Jb�%����d��V�&oӯ���>��}-���[J�b%��b������a�%�z0�W��K��?�d��j���g
]t���&m]����gl<�kc7�qؿ�L�
�i3�+�p%a�<Tσnyy���]ALN��N�1{��z�jܨr\%�rSX�YI�7�jj*Z�:�P��Ҩ{��Z��Οo�c�[�O� ��U�:��W_,,,4+p�~b�M�y����y�y���e�? �^ohh8��D��������酪�4z@�T_��bF��/�f�L�ׁ��G���NVw���@#������_� �;�EE�sJ��W��(��nαӃ������ԘKs���<***��x5F;x����@|��-t7�����05���ʹ��s�����k�Z���{�@�b��'����;Ys����Y�h�o�"�
/�ꢻh�xx��1Mșe��@���{������s'''���>d�(���`�-Ǐ:��	u����vss���p�ɴG<!%��@}ԙ��6WaԽ�``��_X�C[ۼ;9h7iy���)'�?]��p�u�#�r�}Ū?~փ�wf_x>_S��}��.$%�=�BL��D�
���:��h���-��	$ҙ��tz�,�r}�̳擹...!�x%�t����14d�]�E ފF�Z�v-��i�ˇ��?�Мu�0z�┡F��gg��<�ϏB�^���)ڐC�(֌ ���zf�L|�d�3�!n�B�S@!���_8�9�퉤f$%��γ�:�K���ӧ��@��J�jt�]�������΀�1�
��o�j� |Ɓ��S%1?���{�>G��)A'n+c��}7h(T����F28j�����mޫe�#h!0��Lt�!�>Ԓ��o%]�U.<�8���Y�T��3���=nm�|�M�UVV��}�h��*�^��y~p�J�攉�D��.2i����נ��y���Ĳ@z�li����]�Єw��"N0N@�Ǻ���B�y��a!��Ī(�"����0].-˞��X�_m�����]�a�gt�fXPP��n���a���t;�x��S��c�P�.���B4��o�u{�W�{���<�y�ղy��X3�n�x�n[���qz���Z�#A�J{��ށNM��m�))�pU���ХSM�O���g����Qk�J�j��O/:�RD�1Q���t�#�H���ѱ�7T����<ۣ���TG�D��C�#��F)㹢����F���^Fx\usU�����6 �5.;;�_�[5�١D.@��ƺ.�W�������{a&yr�s)��PqԿb��hܱkq�&[��@Y�Õʛ[R�q�G��(*�u��hN1M�	�~�$pjQ�ӄ�����g(բ�o�,������t�:ϩɈKS��@>��>[Z�����
��-��ݼ��|�wrA�^�P%�u4�=(����1А�C�M=��ՎQt;�6�u)���K�X��N�����	�ݑQK����_e�����M@!�6���G��Ί������x.���II4�)��R����GC�l2>�QDfH2�Lvh�R;e�������u���y�:�o�t�繯������B$|R��:!�J���UZ�R|L��_��0R|���]< N=�{ ����?X%����f�R�� +��Z���xgF[_]cB �F�z��/��eΚ��f�D!O<�3B^�s`?��0InP�W���	&��|����Y����&�#��� vv�@ <��pX abK_��~@a�����C��lh8'hM�.�.��������݇&���mg��
C���zn���H�UK>/���ֽ_b��c�W-W�Pj�P
�x3!���BPP�9U�9�I�cs
��A��K7��hvzB:̜(�0g|�Hv���{.o ��yvH>yC�A.wmE�~_�꿛^��L����=�)&�k&� 9~	�+���;Q��Z%xnn�� 7X&e�U0��i��o��.U���^��&:��_�45��;0jb�.�#�m����� ��G�RH��^���|�YX��6z��3�\���+şU���}z��p��x�)�����-�� � Adk��T�q���J�ݗ�̷�h-���"B�A���̀����,�N�c؆��e.�E�J��giE;�ox��@�'$�л9Q�$���5��$���O]4D�@����?ž�"%E���&z���N�\��%G�=A����sߘ�r�K���uTP�����r$C1uj@��5�w�+r[fe%��w��7p�� �_���p$WF��fd����.�-���c�&�(�g� ��8���-t	���/.��d:��CHB��٤����38d�i��Ū�v��$��>EDx�t�ގ9Ӣ)�RpƓ^�eN��alZz,����.�ƺp|ob$;���DK{%�]B��8�E�:	YU�@�ܸ%�a��*X@�dU[�$�!j�Dm0�����L�cG\�?����1�d�jz�Uˎu,�Ȃ��2��Ճ��$u��u�/;^�b;o"�u�핹@�f{�i�.f�ю�۷� 1F&�U49���ѭg��1-�LL��P�JF�V9��@�FGGg�dg������2�YK��fVX�\F~:��ي��+����-���}D��ΐ��ņ�Q��7^��mce=��?;�z|�x�w�Āo��n� ��k6����<��!����9�o޼�(������o�6��y�lXDj	�S�6�\]��lw8v�ko �?E]�W�)������I�?:?���>˹�C�P>�{R�>���O��V��q)��ߍ{{XSS3|]��S��2�>�<��N��_����$ �I��ΐ$Ȯ�n�A���5{�1��:#�m;7�'] �<|�u�I�����"sQ{�-���~�n�Zh4o�q�z߷��߿�mFKU�6�������<A)ybQ�0Roݾ�XpJ�Z��g\��������ׁp�l�>���	��Ouy;�x�``b*�=-�
.��VZ�(�I�9j��Ӓ�0�ݡP�39?^��#؏ǐ�\�A�dP���&�Q5ʕ �~?�e&�[��(��KT�mX�?$�-˯2�����8�
Ѻ�$ݳ�����ҙ�>�^~�o�����Qkv���X�_�� z��.��o�a��r���r,�2��ߗp���c=�9j�؄QYO):I����\ؘ!�q�����F/���r�	����)=z77I��:����7��㄄S���YJ�룑�2���?>:�%��_���y29�Xu�� I*��n���s� �6o��4���*��&?F�k*��c;�m�N�vݻ�T%�����c=�+��3�L���Ғgd�pDf�8�i�o��Ls\�/��r�2|qY'G߱cǏ�������f�e��O�]BPn=�G@aOmJ�P�����V{��e=�M�-dwB�[?�s-�=�jɘ&!@Z��(+W�9�Y��n.���}��"����Z��ݎ�Ȭ8&��4��_x��m�-qII���BB��V8�$9V�����*��&CҴ����z���f�8nyJ��B�s��8�sct��CX3yNG�����r�%�OMO�H�hb���C�4J©����-Q���z����d`n�+2ˠ4���F��$Q�n�U{<����ى�[�wF�d<XV��۷y�N� e`���O�>�:�}bXғ�a��5 <��.kUR	?3CW�АM7��.�𕼛���Fql��B�U.'�8�髫��JV��Ms4vjl;�=����5�L��$>�^�5�����%��I�������.�\;V�%}�{�,l0UO��N�=۷����\��$=�^���eg���o�|�� CF�L��Z�o4��}�LWTH�2�oɁ��m��!�e�$��A��a��Wމ6l�va�7���˅��}���]rf�mƕ �X��#3�H�{�.�KT�?��&f�7 +k����e=#���7�(���S�9	��*�7�r�0Y��!��KM󅰠zTTT^�4���O���C�K�ue��0?K���_{��" &*��]�3ܥ�nt�4�6���?UFI����eӳ�h�U'�w���Y��˗�KMh���Q���;���,3�v�,�s�M��^�B%�R����?B��_���?�"��[���+�_��Ţ�s��)��'g�M���~+K˱��ӿpk���V��?�_�� r�eϞ=Cu�q�h~i��j��w~d	⺶�����mpI͵7�RӑL���?M�dو?+'''�������������[�I�Vs��.�P�yuyyyk\���\��Cx�q�p��%��a�vU�/�C"�6�����ƥw� �f�	 ���F�C��Z��CW�M*Q�Osd���N ��<���C0��gπ�6?� �T\`�V�J���O��|��Yz��b���ׇ�KT#��8��hj���Ϟ�B�m�G�ؔ� �3k��y���z�H��j�Ĵw"$�~��j{�u�aY��f�CV^�ex��w��fh�z�=/8~���c-��o�~ջDSm����[6z���������m۷+.��c�������4����M@91�_�!�d±tuu\��{R�[�����7* ���օ_����m�Bg�ZԡÇ��.%���{{O�ɈM}�bD;�mU�"�ʁ������h��2S� [���o�t�
'N�����08����z�/R�ɝ@�H|����n���v��jt{d/Pʅ��Dy3��*�[轎�k��@޸�޵kW�'�CC)�N�p`��V��~hyti�W�O�}�I-�w���]b��+��P���Է#H~����RY�j�[�?���Y'CܧF���bf���R��o:�����K�����5@��-] _�c��C��1&�x��'�=פ��rT���H��L틋�p= ,���۷��ՁŐ�]����÷z����Ar(���@�Q�j�N��jua6��#n�6n#�T��twJ�?=�Y�6��o�Y��}��v��R��?P��9�n���66����u�-�0_�~��V�(&����p�g_�g�� ]����S���<��e��7��l�\^ªl��ڌ+�O�XX��!�q.6�=`���544,����۷�RRR$%#������b��Ϫ�4���O&GkC!P���寣%��@�f{Ovx��:���1��-,�p���l`ͺr�_7��Ν}�Ϣn���xn��d�;v!8Zbw�2O�._L�sϘ����@�_�z3q���4~���g98�^]]��曟�T4܍��x�p��|�ďP-�p�R�GOx0^Vm�x�Qߩ4��qe��[J�o��@�y)��x�|�""�֍��A���{�qϛu�����Ƞ�?ùE�xFt)Tde�?ߞ�![���$�>�Z �v�Z���A�{d�Rr��/��q��:T��ee��ZHE���3�Q�K����ϟ�;�(,)ImD���NV����&*��,i�E~���v ڏ��ޤ%)��2�'�՝�/^���U{�����g�<������b�_��n�����Գk����=q���Ð
�P�݅�~�`�ܑL`���7������F�&��CƋ}^������]�z����*x�G������e���֢lB�鞧��*�}��vƯ/͵�C$8~l�i@��m�e�@�=��ra��S����.����9�G�j��k�_��<����,��(P(��Sa G�8��ӄ���;i�j�4�*������ֿ��1�v��p���J��»	e�������7̾�_��A�Ha��7?��խ�'qS�d�0��ٳbf�$�[�%����\�R�)�[��2�Nl����gC�V�@x����������?�@?��#Mc�p 䐟��vh�JM�l�PT��|��\aKx��� �P9��(�"�F�+ �����ȕwAk��� �I��"S:)5�u�����:�'>�z���Zp+P	��g��-��
8i�ܟG���m�K��J�#�nC��c��\����w.� J��y=�՜ǏO�5X�6���'��:c�*��*���� @+pL�����~�_;���?*��M�;�g�.�	������mhW�&�#Oq��Z�EԒs�����)��z��ձ�(f���/���d��_�КRo ;�&)�2�v�-��h��@��	Td:�|��`PU�7�/p�"~���^� VNâ��� �:������'Ũ7���%-���W&�v���M$V2q-CO`~�2��HE����6�<hB|��.��/5Fƥ`����K3�f�ZH+�+��WC:R��@�/p�� o'<�����P�u�O�������؁�i�Ro��T^ n������OEK)Z�
�O�A{�4����>J!�%ʳ� ��K������������02���úg��"�U��D-�
L���΢)�+�ӳ�·m3�w�a7p�
����:����􃯦8~� �0Q,�^_�h~��� Kyy�ͧ��50�cWP桰S�s�n�Bs�+�b���W}|�S��4�/���D�_j���|Ll�����6�^j"�yr6B���'n��Z
����G���L<U�θ���L�;���"��r.T<K�-*:�cǎ�dH;n�>��/�;Z�L�/ ��΍������HVϑ��G�%ݵ	{�ΰ	�K���ދ :������0��s/	��� C�T��S�Y�X��!�n����!2^
7p{�o]�(��s���~��(�NC�7�+��R��_N�X
����Zz ѭ��Au;��#LSA�� ����e~�Ǝd�'�������M?������� �ws޼qVו���?�-��p(��վ0��^���p�BNNnW��8J�W�'	c��qp��ơ�(�����	?�	o_���K�8��mI�	d�U&"��pa�0�Gˀ��AzuLN��II>`Ȅ��Ԑ�����&��I;��	��	pX��b/ZH��9>M[��N#�զ]�?��T9����U��-�pq/���ON����ׅ<IKĊ���TW��lh�h˹P�_TYYy���ۣ��?�r��C�i�� Eh}r�2�I���<ذ��i"6�X��m��F�s���5e��9� (��c~�����V0�n�a{⣎���)�����&���{�攼2��㻜W}��!�J?GI��5��?#r�*��v���@�?��W�Z*��=a�V$%.!1���RBOY_����ؓt�Q�z�w��c��˓$�L��d�
��M�})fg���!������t�**��/��=�(v*[��m؈��e�C;7�>�#�U t���2r)�0�E_u�R��V��XV��'|��E�-]����\��!��G����h�ebR��^Mx�쳙G���c}%Z�}��O��}��8��2+>�`82RQ] r��S��r. ��{��Uؖ���3�jl�h�2ݺ��}h���i���x�[��������W���=�cIii��Xx(�hޘz��>��cW�=�O�GՅ ����g��e�N�Nҝ�8�5s�#�<p����#���mL3\<:��`4�5�\&�p<B�ǭ[�rm��r�	d4�eB���GO.��K�;���(�I#����w:0�K0+HZt�%\��?�^�q| ��c�˶' 	/`.����ug321���?7� �bZ�*p:sWWף1��ڔa7 ����!&����6��P;�<g�b)�5`u�����^�hrum-����C[����\��6��7U/#J.B�>z�v�y�n�z��M������딟8+d�ŷԙ,Ѷ}�,18��������m?��?�j
1AW��8�ަ��L�E_�v�Ѩ)B�$nk۝��G+�[5�<�^�K�� ȷ���:F[�ɏB�f��� �LCG!���#�ҏ�#��[e���������7xPCGGW�m��)0�S �8��� ۦʏ�5�����	������%'��/��?rm���o�3��yt�|g��C����Ƙv��`�&�G����>z^����C!`�<�i,�Dx)�d��N'�n������!��K9L��"5���Y�>E7ǣ���QY�J�n�l~Dr����5
lw
���gn�0�`�^�k㿝'
�X���!��֯_�F�2�3z��-�}iO���Ƅ��J/3���B�
���"��@4�A��.p�]6
O���3�%*���2���(G% ��o�J3�.�Mᗤ �P�����a>"����u�;�U �����Te�Gk<D1I�TNY��Z�S�~q�T�7������tE���e����:y��U��c���Ϟ�5e��n��Lu�G�oj���X���
����5Ҋ�̐���,n��O��a9�a����98���6f�6@�������]�r�	8��>k�
ݢɻ�no�K�K�K][=�o�)���wN< ��p� %(��9�Q��?��¦J���qZdhz����@�2��������d,Q1ng,�� �k���)�/���ڵ��X��|TBu�i���B�����NN� �����"}����v,LF�����\����ۯƇ߅�����
5�*~�l�u
!|� q�aa2�͡���_���Ɖf��&��is3�l˯Yݾ���V�rS�/���W�-<�N�4����U��w�?���#{N�����>�c�.���~lFQ�
j�紴����x|�����K�.������;-����gQ4a�?����XPFU��D/A�/]wVo/ ���k���͐GX.������>Z-�&N�' -,~�n�F{�-Xd�CW��S�8�'r�D�-Ŝ��yFSsK��!�F[���t�+���:�y�N6�_���l�	>"k°@T1o��������X�pt������{���UiJ���lP����+��~��_*����x�O\��ć1����?R�b$O~�h�sҌ�'��sH��IX�é�ʩ}C��D�~]�`|F��sá7_��6%�lRr4ync΅���є�٩�q���{ݣ�^{9���:���h��|1 |��ӡ��)�t^��2Z+��auL�K�F,�%�D��3yQ.+~Ϟ=��W{Ym�ܴ�eN���}���A��rw��s{/C{�YCSbN �"zO��Б#���⡡���Di燦�&���c� Inx&��!l5�<���+p<��ק�����~��H;סҭ�g��E���cv�������8m�c{�9MMͤ����t�ܧ����X�y������CG�5�9 H�ğM:�����#A���﮾�~���L�Rz�\���4�|U#��U#�Yxȑ���WUVZ��i�ٖ+�B��1��t��z���]�q�K4 �䆅�?B�̚U�_3.�����su��Y�Ԥ$�S**�	DΡ�������B�s�N6���֎NN���q`!fu�uOO���GK>-/~H�W��`�� A����y�H{;�(+m�h���ڴv=#crj��:?׏�k֗.u� f;5jm�QN�QbX�^C\*L�g�LB���i��7^?�����l/�ѱ{����/�utt4�X�ך�$R��j��p6st� ��8������������[�9ت��-x._�����Qܔ{5v���߽F�R�3�����:i�?0DGGE�������8�ع7ʨt�hU�	���E�=u|G�^X_M�i�Y�ܹ�Q�����S��f��o ���\�����z��	uX��n���ƀ2O#|��A�D��ޡ��q����̙*ܱ���ccc�Wv���ݞ3Wa�1W�^I�+q�[�L�� k�G�Y���0���q�����dc������2>
�Z�6�O�٦R8?;�udWv%�r��I�[�o�<x#Tco<�B}C�����w'�	�9����8cĞ K���J4����s�N�k�
.����/��,$r�E�q�������	���g3##�-[�$'%eTR�G����i@g���-`	�3[90JV�i]'��yN�++�ǋ��qc�3�$��C>7r,��aa3�V0�y�@���} ��ii�v��ky�T�1��W���Ӱ� (�ɱ��\v���*�m�--)M*��LNJ���۰���@ȇ_��%R���wr2����X������#��L-,
w�<��D�%z��L+g���j¬R�P�� �eZ��>� �댾~
D؇	�^��hL��Y�<FK� 듊�.]����]e^ �Ԙ��}�)+�k�[y�T^Q�'�N��t2P��`@/�����~˶TwqɃ$�TRR:t�h���OUUϊ�ǵ45C��#���z�8Kz|_M��/>uY��l���ZK8"ki?�H5Cô�EuM� Drr�ɦ���22P�����ej�������v���F�\5V[Cm�+�Y���Cx%����}��b�Ձ!��|�������k%Jnl۾���s�(=��ZM������b#��Q��rj^ޟ��"�: �C���Ϣmu y�#�=a5v���yᤦi� "��˗���F��܇�œo�Zm�x�t�Q No!��V?�]��� J�X|ݿL�Z+�}aEEJ<��Ȼ��O ?L���j�N�۵\�J��Aܦ�O $?~�{�*?˷�x(/����7(9������u�#62���+�	iH�5�"�^���.n�|�a�G���Q��Tյ�,�R����c�PA�z��H�'c����r T�����2��Pd�-B��6W�}���
6�m��66j+n���.ζ��=�ho�]F�l<5,��v�����)���B����㿀��Q��c*u^��b!;H��7��T%X�L����S�<�W�D���ˏ#�ŖVVָ7��oO����B������=�~�~�r%$�Kh��y����!�N:t�p�uӎPy/N˫a��6��d��mx�P{K��t�j�����%u^yS�N֩'�^�^��f���$��g� ���^������惨(x8}}l||��λrZ:��VʪPѫ�U�G���i�K1����"|%�544���i�����n|@D$^���DH�̱a��W�E��c��2^�ƌ^�g���+>D?+p��.����+W�������?�L�:(-���}�*H/3�'K�p�L��L��7�{zzL�)�VB�p�Nj|}�NDJ�r�����S�o��ٻ��J"̏�����BV��ܭ��wfh?�$��PӾ�@E��d�TE���x�Õo޼)���~Mw�2��J�vU��а]Fզ�@rW��'!/
'A���CL�$��4��N���[�!Lm;�Hg���������t�ۡ'K;�^zq~%�)�k�����=��gf�Ё^�ƭm�֬���M`������Ǐ�����'���y�Y`�.I}�]��n1خe���U��x�����f��bb_�|{�X>��J[,|�_qH�y�l� ���I񨆠=���l]zE���4���gϝ{
��e(Q�?ZRB����x3�6ˡ���� �,F*�S>iz�]��(��6m(�A
�/_jn޼y/&[5'>x���0����)������#�#�!0uɐU7O�:�������/�4�?RĦ�I�/k�)&(�����i��>�Y��?���

�T���$�yxR ����i���<T^�{�����`��E�÷�gF]�k�@����SI��
�qEE��g���ZO򴙛q�D�DA��#�G~��i�����(`�+'�9�o�n�6�P���&
G������n���f���1� -���`#n�x�rhjc�Bf���k��}��}߸�+��0�l��g������%�~�U��NR�䴓����ۇ$$@0�U4����B�^�9�jneպiͪ"���|�r'(I�|6�;�G��6�zW���VffJt���}��R�d�Y��"��)'�j7
���ب����a]� l��T�lZ����%����+*Є����_��i�\x�	lX3#��G�
�l9�l�����%�m�Z�;��n ��`��>*Y)�k��z��p�����ϩYnV��7@�N#���c��4y�T��7�\�aq�0�����5�rE�F��[�����L&o��u�]M�r�?R�����X)e�/i���r��1����@X��O8�lγ�<0 ��J��gm�s�q���AѬk�F�QsO☠��������� &&g��<�@�żf�l�~���/[��z��*��&�)����߸�������[xϿ<d��]}c�|��tL:#�pK���-e].�+��l|K����<ad��(l
���m����~�E+Aj�o
)tJ+O��edo�:ꮓ����kq��wJ��)�I�ek�KZ>xP쐘��Z{����R�Bi<h�[|���c>M�I49)6�j��ݾ�ٚ+%����3�*`"��f��ϭ@Ҿ�S����y$��;�S�g ��@�/d^�o�MD�>{�J����0�g>�YA$���� ɮ�M�ku���07�jXl�\mN��Ơ�C����xJV�K�&�V��Y3Y4�g)C��Հ=�]�O7(X)'n3����@ȝ�o��ǝ��ux+�u�h�t�}����IJ�	�;�<�>�IUM��)�������Fh��e/��J�׺x6��P�d�U�a���m�L9	ݙlj��s0�u���'��ؾ{�g��-E;O�]�Z�A-��_�>�T����8m9�����oJ78Y�rXG�0�2AwJ�롔jՈ��N+S��⊃��S甍��v޳gp�������>���=OZ�wԔ��M?�͏K@�������Y/�`�6�|~��Gޗ�9 � :����&"N.��k��v�>*���Z%''W�+r:�(�2Z���d�߷�@c������ni��_���`�O���|�T�� T�
�?�4�q�pkk�����,�\+K�_�⾊�`i�o�v����v�[�i��,�D���}r�>�_��@S���-�F�y5�%<|b��2E�9�F!	R<��Y;������$�{ |��ׯ_���D?��N����#�̷;�.��f~�Է|�U��)usl���sz�P�#�p��]$�C���QD�d4OI͐�!��躈�&@(�Xl*��v��(|M���\���\đĪ\�G�8�����+[���{	W[�_R#�9W�-�V���L�;��R,���H�#����Bd���:���� �2V��UP�w��5F��|X�
"U�>��γXE�%1d���BBe}�w�"n�+@`Y�*���:\��l߱�,('
���vDN�.r�>�����Afzb m���41����ϡ��&��..4�'��^���Z*#s{{KKK=������E/dhG �0��B�����t?&f>8nB��2H�2֎��KF`/���ݪ�����PTDa���o4y6�Ӥ���[,���s��I�q"�<]Я��m�i�N \\h�UY�*��1ӟ'Cċ8䐅��?�W:�	Z�\��=ga����R����!F�%19�FY�U\��k �x�U�ݕ�=��H���{(�O��\r��_/-��sp�����l�"T�>\���g�$�vs�7,j��d�Evܝ����7F+��RG \��|��PPD���/5�_Dt�Ta��7��_���.N��bs�b��S]�e6��87�|)LSދ�!�1�+`Pxem�9���DFf�w��j�;:H%5��Ё5�S����e�kf�y�2�m����=`�]�����MV���^�)WDB�V��^̲#��hg��s?��h3��_���ƻ�?q�T^�������3���,�C�GG�V�@&��۰�JE�~33���̙�Tw�7'i��.J!�!����ꚓP���K;�� ���_�}s��*�l�����t�T��h蟷�}�8 �������X5r�����s�`+x?J�R�V���Ҳ���X\�h�U%�A+����A��yq��cs�U�	�ϝ۷���]C����7�������@"uv�P}#���k�@�P���{]F桨uC��7fz��v�L�'���&B&�х�閝�>e0�Py�bF�!�NPP����jj��+�~�a�"w-���KY�A8����Q�����b[D�����=��:�h�y�|�H�+�ʨ��{�c��>��&�(�bee0	���z��yy+u��Q]}�L$C��B�gY~;Li�Nܿ#��A\��>���S��L1M1��5�,�����T�� ��ּ%�ɉ����J�~� vɽƤ0���4�%o��@�O�]��&���m�}�iw�8����z�*W�}Ce����.���b���zl����(2[m^��v�o�&n�jJ�
8�qF����5ck�ĉ����2_?Ŷ�.b��D�;�nD�X�qjҮ-�D�j�i�P��|9ee���̳ccc�II*ܱ���!�z����ف�LR��HF��ouu���v�ͧ%��Ƴ/�Ӹ6P�ïa��>��-�i���Լ4o��,`~.� %J�ɬ�c(D���i����b@l��.��}(Hd����r49"�c��� �h���+�'��bV+U/C���xz�!�@hX��ݱ��bf��L����!D������t,~��VT�- ��%$(�sqe�2�脹9��~��n2H��ݻw��:�_><сv��t%?��V�����*�hd�����hPD�J������X���6e�&��_��d��}%��kw|x�m���r/�Q�MI�וB��ݴyXr�<8�P^*�2`���K���gۅ?u��f��X��-Ƃu[*��]��H���L�V����к�����_�+�]~�4ɪZ0����N�6-O�b�����wRJ�ȡC3[�H���#~@sr�����k��������[-φ=�: �����2����כ�~ONM�V�
�hm���K@���G��ސ �ݑ�	��<H�����QK|�ܮ1U����q�ӖH9���Lk���gF(-���v���"�{R�D0�؄ːCs!�����2,.*s���/�I		EQu�#Z�韖��a��30m�j���G��W4A
_���(���z�����+��6.!A��	���_��?*;�N'�85�
��K��P�
���p�`����8@��cO߫�݆�KH���q%��m�6�92�mX�?�n �����uO�6!����\�y��\�5���bo�R�<�����[�n�Eu߾}��}�^^��>ѹ���$�Կ��,F�;6�R�0���QҞ���P+���OC��3�#Q����?��mB<=���*�x��p ��ڻw�9�$d^��.4X�ҏ`�v�mK��S��Ptv}gh�*��@�PGd��;G��J��{'N'C�<.#cHVr�IA(�A���.tn���sUb�x������}#N��lR�R�����_]^Dv̈븁�����w5�~*���A��y���:���Y.�%�l�6Z� �_5��x ��\�	�����^@\槗����.FA�쓣�����4ꂔ�nv%�R�������y��ˣ����(�������7C�o�N�V8�>����Gi�J��T�[:� �oq�����III5l/	޻�i���O3��*Y5mK���j�P���k�zh.�F"���M��1M��4Ɂަ �avʡ����s��J���7�xA�b�Ix���&&�1k6P���G�����HN&:+Ҳ�ص&�ҠM���J�#"#5$w�cӨ$�K��7����c�g&J{�k�o�$ߜ!y|�]������
�S��[6d�9��݀ ]b���f�H4��`��E���[��G�II$�o+�V�^����GZ.��jr8��7u--�WV��41IpXmS������u*<�H��K8�k�8qJK��9������p���	�
B>�i��D���е��%��EV��}���A����<?H:9Q�'���V5<>�'f�8���3�:�C�8�����	��ed�%���d�=
���C������)�	 �}g��fx�?r#f�q��|�N)���S�������N�� &FKh��Fm�κ�hh~N~�T�/0Q�RE�f��Ν;��w\�J�&&�̤9�ʡ��78�����^9�K�������k:6�vmt�v׏�6�鑨��`��K�&a���ZS��C���P�N5�U������������D�[(a������T�9�G����_�~�����nm9�TVx���nAV���w.E ��Pl�#��n!
�y7�qKA�
 �� ^ǼT#��zI���|��0آ��ޯ�ꚰ��3 S)zy58���˫��;�j1�!=j�l��̰:��ePp�MITl�	�}�ݥ[݆|o3���-B4�P���(-n�_2�.�}9c?Z�,m���`��M{�oA�PZ�T�y�����1��ގH""��@�v%]���%�V.�ln�۔���Pu>(*:%�R���i�H9y��_���Ygggů��p2�R����Қm;�t~��.��D�~�ͱ:U�1t"���'c�CGŮzq�A�;�L^]���p�=;UPw|$NSG�sօC�2��;��RH|��xWW��l�
�H�'��Y���l�ʪt���޲�h���?
Tp7�sݼy���g�;�XB1^���+jx�N'���#<+Q'E
II�<x�#�޽��6ɪ�W}K� �Aj�� +��Ӑbl+��[��^:K5f�!�p`��ñ�n����཈�9K
T���ym������o<|�B�X���TV�~�e�~ଢ�"'�7].��G�Zi�&2Ujrb�)���������	M>�3y�O��|~�����R�?z%�;H~w����Q�2�����xԹ�5�
�C����.Ƒ��ٷ>�w�+��c���N4���b�ݿ�/�	�z�ŋe��w}_��2gr�T�%M��s���km��~�����Ѭ��I��_�͕JM�9�?�3�ƭdm?a�3H�3Fy��+\��CV>�Cd��,��R.��*�(�:;ָ0ә�^_W�ש?Ov��q�q �:�J�D�-pE��jgA�/[mi���:��_@��mג��
�̾]��	���:��	
�m��􃈈3��)�v�3��M����b�Dl" �Z����A�����Z����z�}�Ē����/I^��s�ކu�����ZZ�6U�](�*�vqg����y�����;���=���ӞϞ�7��&l�gW�^���T,��B�y')���˗����z��h�ꩱ�-�&N���[{:?��DoU�JP���
0|˖-��h�563��q��~��`�n!��V���ر}��=m�Y��m�O~ ���d��搐l2b;����۶��q��Ya}[[Z^^���g��{?W���l�ii��.�O��ZC��)$��3�¥fn�k)�jI�?���ӧ+��Ǚ�F���࣮7kۏ�)J��x���Wݢ��#Em��>^�������(�y�@��S��gׯ|k�B{��s����������_��6��X�YJ��_󌌌$'%��5>]���eT�6��Lb�S^�������<�3;=��=����¾5���Bu\����MM�&�o6��'�1�CU �nM ���������A�13'P�w*�\/)˶j�*u�����+�&)�j..D9�L n ���M����
=���'&5XBI���{57ջp�F_YWw/L�0U�׸��	����~��&X���%�@cq�x��D�D� l����z��A�� pd��17R��܌�˜(�̝>f[�f�('0j�@����2�~���"�@tUwvvr�S��wǟ8Z*NM�R�dl�̓{wf�k���/:K��.xJE�
�T������*#�~��)=Upo��a�/�*�g�ޑ��,����TFI}W��l(+ �Z��?	Zн�yͪ��jBˣ�F�K��b	��3�ZGv�ޜ9�{����mƖ������90���AV���Q�[(�[����*�&2Rts�@�?C�+����ݸf�Ax�:O=Aua�kɐ7�B�~},E��\||��<m���p�$gq򒫫�mz��N3RM��Y/}� ��`�i�Y����{�v{�Vғ���M
�!�!u�7���&f�(1� �Zq2DL�0��G������Υ����M���K��M}?D�Ĝ[}��g�L�x��έw�mD�9�'�mx����[4��rVlJ���TrJJ}楊�vF�Q�x���O�L��P=k�>�O]���[��lzA8B���>�o��팏~���c�ž�Y�&�0x=s"lcv�L:{�r>z����jp��y��T�*�������m�!z��#�ǁ�k��YHo�����P`XA�>Fȏ��w���'GN�̟��+�@<2Wu��/�_�ǔ���V�^=��p���~t4+��3M�ƶ��	�*�Pe˰��q �"��/T���%!!�c�4�� ��*����ٻq�)��9���_�Q?-=�9j%j^ Wɉ�镯9�$O������������{�Jrr �{�|����cF�C�$��/E�߲���/B��	�Щ����3�m�@g�������<�A^JŒ733���������Q ֊�2�ɜ��)`D��?��� ��voӂ�**~��Z�D8��L���t�\\x38}Ba*gik{������H�N݁�����	�2�wEQ8C;#�SZj*MM͖��*+?N�c��:|��8p�l�_�.�:��)Ο�C�$����~����ͼ����IB9�����P�)�#�n��[Arkhj:&�',|�1�\u�巢��������D�9�}z<e�*j���"��ϟا�\Y�<PF�jC� �'������W���y)S}���v�Z��K.*2���ZR�� 3���σ1� �K� ��?���l��8�[�'��Rr�;䌹���7������ۗ�vNQ��\���������Ӿ��u�D.p��P�&ƾ>\U�Ԁ�5
<�B:������Yr��Vm��j����։���ӽ�%g�����9��d���:i�F����R��}��"�����.I�>�>}�܎�)E���`�1]�F��i�y,�E�oY�%zr[n�N�cwJ���%�~��|�m����1����& %�I��\hhh_ ^��(����@h�������m�tC��ԩ�fff,�D�jɶ	�?�Z�����+l�Z.]�U�k�LC�uOu����X� b").Nj��zxd�����tnx��L�>���x��:|��SP��� 2�Q_7��n�b�X;n��/�t�˦G���ǩ�������%>��SΛOK������߿g��v�6����C.U�uW˳�ڭ;�p��	B���nb���+��9'^��#�5:3R5���D�A�\��! G�4o�����a��}��E��>�y(�E#��UU��u�-��� ����ɍFK���ԇ��'���&0��ܐ ���#k�X9��T\l�����#]�?33S�#�������(�T�%1�h�����|�׻ncHNMU�n�>1x�c�.f�9<ea��ʆ'տ.+��i�O
���oV1[YJ%]�8.��c�ܕڧ�t���T[?\η�ƹ
���E�qnc0��w�~��2�J��d�������V�b��{�>K+r�y�~�IuP��Ҹ$�;p4���KK����5�x� ŰӸALQ�,�y�	�&FҮ-��_��v�XN��g`y�C��.P���Ggf�jcf�b>��%�kt���xAp�x��	b 1���G����?ĭ��+�{ ����(�F�Cބ�6	�M�u2��	�Ò��l��ʵ��SJ����v��h:������@�?������JUn�j(N��˧IGFq����1l��r���y�\�k:��LRq�%����N�~�
+׉'���Vf�N����\�T�S���i=-�Ҋ���L�}��D�$cg
���Y�G�&�ɧM�pqe�eɹ� �H����9q�&\���vv�a[�ȼ1���MP ݄�����Ƌ/�u�1>�����5ӿ!I/ �n�g�+p��콗U�O�|���58�
�&���//�Q���,;������!;v��/��#"��r�xP =��;�A�}�����9��~�Õ�#3d���C�g�3��<��P�^����=m��'T��'cҪ>J�N��V��x����]�kX�z��sSc��t��akgY�1�p��0�;q�g�}'4ybL�m��)��/6���e��c;�z�$��[g���;�-<��>U����9ǘ��%��l�6+�h�]򬬬��T&^-p��o)�Lk|�e�9�"d�Y��[���E��C����ޑ�_Y4�� ��30$fg;V|������4�7��8	�.�����\U�ٽ�pְ��K��}2�k�Ξ��c�r8�ӅeRKtR��)p>mz�^bz��wm//�agIeWG~�ZZO�1���ފJ��n"�1V87�Ϝ.�w �W7:Z��O�e%y��������s鼧 �Q>����L�utlnF+ϗ�J�����_E�۔�?m"�������k��u�;��2 nB%�o�1��.���2<57N��s��-r������^?~C=��4KS�o��5]]]�� �KI�K��Sg8C����ۯ3z%�4�_0�`�^�>�J��1�ڔ������;�����/���b�H.� ���%"EP��T)"�^�%J�) *b�Ho�4)���(H�EAi�A��7s�����'O���{�̼��̙c�������O�����*!j��/�t	� L���D���IIH<Y��c������%~qqq�asu\�&5���k9�1#�Dşt���;""�q�����O\��͝�]��/
�/��rz�s��`���<�o��׭*5��spYo�Z��EX�̕V���<B�y�!�V�4_�R��=�g�P�߷��,��~�̙�Ç�z�M��\�n�oln���� ���Q+����ꗰū�%��B���-�������}�|@����Px���W%�Ꭲ�����9+'�#�zӋ��KD������B��wb�Flz7��g~�
u--�x��|�_�]@nW����������ĥ�Vڒv�%�wEc
KH����s��ԕ@ >BH����7	����=r�eX�x�L����b�Y�vyO����
�W����cc����
/��xsz�y����}�����Td��Ъ^���u7��prrZ�Sγ��Q*�><�X��}{��DVZP~���c����&�4�2��T��}+U�� >߯�:�-%'G�;K\�>�5dr�R���D�p�s��-��A6>��م��յ��/����,7ۼy�Ӈ�j�d*��"�w���Z[��￿�Ţef&�xš���4
�����Ȯ]����Ľ�h�#G��	�yI�e�/oH�D��{�"��&ܟ.<��KD�?t(ٽ�S)Q������t����<=y�'��aX�P_;��\�U<U���@

z"�
�qe�`�dd���wK!U���H�n��84/-��Ç��D�L=��+c�y���8��{'�0g�޷����		k??���1�<���ҭ�;nCZ��J����Y���E��`SYVB��9L,z_�b\?�Pme�B:��3���ӿLy?��^~i*���Uﻛ��t緾�<3�e�~��3�6���P�vV�&��Tc�5mCCJIgL���<~��]<���"��l�*W7� ����Zb�1t�+�k�f���;������⋗��7�jZ[�]d��.'����:!�'F�L=Y#p�k��;j�yx�}A�?������D�I�7"�,$A�m�����(��Og�qF�'�O)A|�Z[ ��Y���.�Bv�Q���m�x}��� ���>��� �}��P녝"Ԁ�:.1��� �Вx�Pw�A�=�����u`���3ڽ㌜���N�3�lR��I��x�c#�hE����a1�κv1�ʑ�rF)X0G�>��=<
��P����������Ӓ;:��j���&�Z�^�8��[J�������˔�<l`:��=�ۇ�!�j�7@Һ���Y@��i����R���^�`��it��KJ�1��!鏏�Dԋ��*Xθ3��oҘn"͜�J���0T���mˢ��W�w�6͌P*�,�9ٯ�	�ҾL�Nj�����/���(�x�p����K��~[�`�6� ���W�>��h�h4�o�����L@0e�_�7����z�09ӎw�{ttt,��Td���V��Dĭ;���� �C� AYN/r��eV�k�U-�w�Q���*�v�gw�h�o4�[4��x_����f}�=��g��_}y-x�����]����b��H������#m<�B����~�E,�rI��xh��{_��?���"�?!��o���`jn�� ��k��~s�+w[*���?�G��8]��bׯW�,�k���ʅ�6��e��>�O/�ȥA��Z��?���f�ׂ�P8z��o���<LN�%#ݢ�";����c`��N��9x8�k1�盺�M�
 ��^�����e�.���ֲC��w�d��NC�{�a�ґ�xs��¾o��������|������?x�:MϭW����1�$�߭缦ml,L��)����Z�iN_lsᠶa��>�b�^�J�=��	��W�{�h�8��Z�lcN���={���///h�WK]DF7MK���B-)Y����޽{f�`�������P�=�zqaa�~��]a����t~ώYHitYAmC"���d����}jj�m������6oڴ��6`� !G�qvμy�|��hտ�5B�'Ѱ�y����k��p������׻� N�&&�?ǵn�#gᱩx���� ���/�㔡*oi�&AAy}޲!�SfuD��?^v�z�%��U�~�����I���ѩ�]�!v�k�ΝR�SЧ��(\�$�5�{�7��,��;���;�p����Ȋ�1ʜ/C����Ғp?�������׀�/���)\,y�8�o���ɗ���� �����*�v.=`q��c�0}߾��luu1;*X�ANś?�Χ�G�ȘEX���D��L��}z��!kHXÐJ��W��(�iFnO�������Qe�!+f���*y���s�r����qqq\lu��?�JJ8|Ѓ���mmlT���[��Ȟ=:ZZM���N�
b4n�o�A�G��$���)�q��ŸU�%���0��U���~�E+�f`������@^�Zw��?95�R��[C��������[��l�T�`���e߾L'5���'��LZ����l�s�^"JN�}�oĥU|m,�$`�W��Bd�1�P7��1A�Z�~Ud�^]O�|����%������W��X���#��g,�B�577W�q;~��`0��7o��YX�[{�|� f8��sr�Dk��8 ��RU� V�*�"Ew��<4r�ť�I�L�6�R��$t����xahii)"*����#�/G,u5�mkg�V}Q����y6�p�hܩ
)tqan*+%�ϯ���?� c q�0��1��! xG�\!|� wq��M����݇�	�HI1�״t����m�����x�Z�u��p�AB"+c���[X������NW"�Ù#�ɆN!���-�� f�ѕ9�������y�*W�뭡:^�u"+(��JLp�{��l���|c'w���ҝ< R��-��ze��-<kq?|�6e�6�95Y�ʲ�2P�X�9�
p��9~̈́��ղ�։��X�e��tvw"85.�˦FW����O�U�Q�Vc�ì�V4��_�a����_	.7���4�/z7�}� }E�>����j��f���;-����*o9A��]�6��Q�����K_�;>�`5��� �� ��b3,V�V�TwtZKR!2���*��	���8x���B# ��`��o>��2~@��"����
�]�y�w�t���;��/��D��׉َ_ ��ZhZU=�d"W��X=)-�,.���=����W<�IQ=y~`Lz3�QQQ\/�ps��n��+�>3˼;7?�cS/����Jݛ������~iH�zŐ��r���:S7�5�L�z�|���6�q^�4�8^�9o:�N~�=6�>ҁ�.��&f_? !�\�]bco��
��Ī�vl�u�ޝO����k�hT�|��a&����vu�ya,&���!>�7�Z(�7&��O|�������K��i��3�)|+arͲ����On=W>�N��m��.P�2!.����λ���.��f^`��9cϛ�66�� ����oRD�'��><ҹ�ќV���dT�.�oNP��9q�2�d'�!���pdԝ8q�TV�,��g�`Z�h��RRRI��:��G/'<�`*q'md��98P�[�zZM�c�~.�ccImK�܈��gq?z8�xl�̈
'p�y���	���$���r���!����ݴ;���� H�!)]�r������3�b���q4< s.��\��?-������]eq'�1B��Н+�[l
������Ԛ��;L]�P��'��؝T"��k^d井�E޺��F|�t�^������0wr!����#�5��� ���@ �e�4��!Z*+ՙ�eZ\<��� V�W�J�%�W]]]!�nz
Jq5�E'����m���O�9d���Pk���^sS"+�R��iu߈�U�AY�3y���[f��'(mUlOP��}���!���kg�s�M	LX�BZ��������wj'�n�Y{�T��{H��w綴��#z/x�p�F���O�{��H�!�J�Z�E����l���䲎�RSS�hj�6�z����%;�������Z�	Л����������WOh}�t�RL������n����@j��e�2$N�:���`��HV���u-$�Q�й���R�5�R$�7��l��\��;��;\�ߋ��b2Dխ<��_ޅ�:6Fʢ<ܼ��lٲţ�u0��i���ܶK��^͞�B� .|�����",����^3���W	�_�]3q!/-�6A��ã��q)�����b<�q�&'{q�����o��ޠ�|���H��>KL���fE�Fnr6r�l`��c��;�2sT0���,O��0�8s)Y�;dom-��OX�����0}{'<<�Ek�c�d��i��p4=]�ߥ�	���)-���#��%�R r�	���S��.
�������u�����LZ9� mh���I>��
 �����]p��\k��0i����, >�@���-�M�+��0���f��5�ͩ�3�ж���Ғu���4$�''=��s��XXo*~Qv%p��?�z`@SW7(T?�g���Pg��_I'�/�N�hjj�o�1�b����JC��-)�]�y�%9O��}�*`JX<Ԓ�Ō#�b�A���R����&1�TY[G�z���B��ƅy ��J��_�\�U/���Hxb+��{W�h���H����4-���e�v!Z`Y�&�\\
��6�}�u`x��?�����Ȼ�s"�� ��X�W���o��I�ZQ"�cOA�hm��U0�\�7L��^SI����&�
6�lj�=)[T<��{r u�\Us��
1�_�þ��{�Uy�I������m� @��2�Ko�U�-��eU�6�<����6z��t��8�	3���*؃�3��j&ʻxj���V��j5:��!��'g)���*<�x�ȹ�r�������i��O |��OցAH�60	A�y�;�Ȥts�sKR�\aA�ONVbM�jj o`�������Y��Y��0Q�=�$�x�� N��>�2���w2=�������@�7Un-��;��3�*?
*����}��?�t��8<���^%A�P.L+�o�uYAd����p�.��E���3mp�}�d���Cf�:(��mL�O�Iт>�2�a�v��p_:���O;�EY=<ci�I9d�++�?z�pM�]"��>�����'�H|���������N�Xl�|������i��;��9��x}}}s��D�_=�n����e�:oO*@�0��k�"��+��,}k�ゔ0����8&�`��sE^9�&�ׯ���彇s�o���ގ~=�QdK^�"�~�D�,�	:a!Jw~��X<�u7��]g8C����(��/��xpMd���n��8S� e������")��x�����Ek����R�1U��5e3ԔYIN��.����1?,�k����M���������ԅ��L�>�˗/OJO�57
�`ɜ�����iF�ב�		xJ�?ށr{\��$�l����d���,@m/�QV�e�yl�Ϙ2�3�u�CY@@`�ƍ⤂2��-*Z}5�s�vY]��7.���JJJ�-����-.�(�IzZ<��1	�40���5����A�_����51+84�8cdd�5�L:Qq��9'�͛�uu�u�n��YnV �R~��mjr2�y�jee��C!�ލ�0&�������%v�������ZHUv$6b�p��3��n�l80낺KLT�d�E��6����š΁k���o��uF���)�TH(����r@^Z�� ����X��ـ� }��}a�^��
�>F~5����A��4y>���`��gӋ0��W9����W�5u�
³�f$�U�]P֒q�����Ӏ��M���m�GJ�!�V��I����,3������K��{�\c��Bt�(�^�mt�䠤^�5%R6Ą藦�bC�׷��~�]�ڶ��=ǲ�׾9�w��Ѳ5�US����aH�Zi������蚨[���#=,F�1�g����}֥l����h˿̔3_�`�����(�y�ׯ��Ƕ�-!vCǥ���U�*s궶���z� ���g�0-w[����`���*	�̼j�'��ǹ�A�ը��߇�4����K����o��|���r .�X����0�3rE�zv�ER���k��r����+�L���6͌����������f3� G<�~��D��9�
� 4�o�eb^�b�p{�TN��Kk3��$�ep���#:6�G��<6QS~�_��o��.�,�_������k{���7�{�N��Әa�鴱qZ|����7R� 2���>���@�2��v��p��G�;���R�z�c��hҁLˎ�=��D����;
��O�������%^{0��iϐk�tP�F������^L5�B�R�QӨ��N,�!���'�3��3��0NG����8����G��J��mj��fT*�׽(���ŀCh*+ߠ9v: �˧��p.��p�n��_WS�U��nrS���\���ٶ1]x�0 a��Z�-$Ұ�|>�'\%
ӆ"����m��r����j��i�#�i��W0W��{B�f	o�u�:B	���w�t�,��Xl�E���ܹ��ە�_w;c�4�� C`c�Jf�&>g�]�׎>U�}�qZw�x�n�n z8tu��G�M�)���%i�v��	33?���*:�)�0��;��]\�����_\�rYU�V���AeB~�ɫq�5���<�tBۣ���'������h|$(XD僃�]O�[��A������GN���L/����C[�c,7LOяc�/ ~��FH޸	���� �p��i� c-�)��ի�����:KEx3���x��(D�2h�u�p���&�v��w��8�!�39�^�o�,�� ��J�wrss���_��Q����ܺ��
��]�Wꭌ��L�_�2��'�;�}�*݋�"!��u�Q�ub~+������`�S������� 7�p= SO�"�LW�;�+���jg�":��]�2���Ѵ����ʃ_���6y���IHZx��f` ����[��Q-�&�>� s><�-���5>��{n�����}+�QN����p��������)o�Ǐ!���g.g�i���I�I]�/��e���D�ՠ:��dP�� l0*<�ڐ�o��8�)�r������I4�3=�iqɸFa_;�Y�R_I��LC����⥅[�yP摖��0x�~?r�
�p�ӹ!x.�ب\�|s����Q!;����ύ�:�tX���ʪ���X��wY�('�6h��}%cSPw_�{Gu_�3�.�v�!F�ں�"�t���5_*"����/�[��r����Q�/��zz��U��
�RS���y��L����ow�;�cH)&����'�~�I9�8�9Y��OIii�U�� X���\�uMy�hj>��\�2Y�1��������'��YZi�w&W+��o$��\J%�kjƓ���|p���ϰVBH�ٷ����v�3?
1< ��0���.E�N��8Q�P�^��buE��!�oMU 6.r��ڂ5����y���R"`.M�#q;Ò���; Ǿ� �r�����(!=��4z�q�?�r3�B��X�����_/ �q�3Xp���e���E��r����*�_�2߾Y���

��ռ�Ňt����ɓ������MT��c.xa�`��>.���\_8R�\S��jR�tR33V!l�fOp5$˯[bd��;��>�-Bd
9z�	ڷ�)t9�2��%yBI	��m�<�\p�k�!q�	����`2Q,X�W!�������*G��|����!+�ի�A��\���ǟ�λ!{i����Ѹu7��$?�[ekf�����u]���>}�7ҏ O�<k��������	��'@t}B9꿵7�ۍr3���������4�����ܒ����w�S�r"o6ֿߓs�W�mo�>xpH9��� ���/O�������:?h���,�`����R@o.���vÑ�ӎ����H����k��Nqmm2?����]�k�c��4�#����3������ظJa�%p��5?m����uɾ��4�;�-��_�#��w�(T��!���bz� ��:~rU����}���c�̻�>j[C?��
[��880\F�Ŷ������jj��\������_�Z~i���S!��
M#�h��	���I�����R�ewIg:�2p�)`f&��ׯ���9?�(5'�ӡ'��9�"n��ɤ�i�d�������M�~����e=B.(�/,�����-�����a<E�F�F}�YO��斔���;��W�O�>��
{�h��X�}�[�M|��u?Z�щ#��
��r�ac�5X�+m��w<�|�-�;&(l�tz��4�����O�����������'��z�v�T$B� ��i&у���R�T� f����E�������,��8+��Z�J����<vzF\��s��o����0ǜe؆P"���wJEXU��WK$���W!=������..��Nd�`h��b,ڟ$�A�� O�a�de=�=?WRQ��j��H�}�1���%�>`��Ƕ�p��\$/uۡU����(ϊ?�CN��05\8"ц~.�ʬ�>�x�&�%����wmœ���S

O������~[y�������ɝ
���6t@�E7;�(2G�dP�%��LO��j9rT��G,���h�s .' � �|Ɓ�ѐ����.����ky���RߨM�=X 2�4���п�'>�ϟ���Dǭk���������%�|L4��yM�MNMa{s&ʥ`I���١�U�:��H�ر�Rƾ���۸'5X������K�-'�ix��q������zX1�9�r�>�(H�e߾� ��;3kI�����+X��%K��#�j�q�U`,�6�[!(?}:���
��	�2$��ݡ'/���17
z=&l�>::z�-����p^ϡ�F�r�Я��v\�v�Ⱥ܁��||bR�
d����,bI(�d����^IR���O0}�2v�v/�Saf�Nݗ��#8ՖOgXB���N��Obo�P˝��[�ENg�:^/�7g0~�!�D��J�^��JJ���b����s�Ć�ـ쇧괮'=�����>���V�J��*��m/t�>9��#��t�w�(5�2SW��P��჈��\�"�T![��kb�}�(������]�S/b{Ig�S�0H����$ȱ��G�l�eE(�j�%O�n�S@�^=��Y�ֹva�S����'M3�"��U��4��K"�O�9����vvvv{�ln�?����H&�g7�������@�K
��B�%,�k��P�ݽ����YE�G�==���9,͢H�ߏ2ױ�!JҪ����i��*���&�[%�v�~�,6�|�Კ��'rRR�$�g���= �!#�Ν�S�q���{�O���N���
?����㈃Dvﮎ?u��t+8�tg=(��d��DTdѺ��]Yj	,���ߚ/fgO<��E(fl!��38�ּ�F�o�KԺd��b������f��$�l��r������&Է���r���J�&���݃M�S����Тo�Z;F��9�:{s�0���܎~}��n�����aq�s�;�ը���3F��J*�du�=��������,J��o���X����'>�#:��{E~Z�����z�6�cH=R,�,ءe�5��@6uO��b���t2r&rlI9�'���� ����Gy�b�B��P#��u���K�-�ߚ2o����65-�~�TT}q�H��T.l���$��jq\藏@���Rp	�S1��#8UWu^Z2dCY���{��3�iU�U4\�^���;�!�r�lT�����т7����άL�$:ɤ�<�o0��7�Ly1!\��է�m47�W����ց�Y�����Q����-��]Z�.lE!Ўϝ����蜍��WOHW����^�a���w�j��2}��ꑡ�|-��8o賦Q�'��[==�y����ׯ_��m�ul�(�^���0�ai/��M/��"#è�m!1���Qpr�4lt~���;�wtggb4�>�+��]�����1�SSz&f�+(�k�lWƭwSй\�,�c򍮍�nn�Q�<�H����hN^uoo��=7rPg@l��L�G�`�'/x��M.,�k>��\�f������gZ��R�PM
��Ɨ�+^������Q~z��S{�r��~���^_��HYI���|��4ly�� T��nP��]>}�)L1~��'	³/h�@��$��WG��=�6Td���0ľ���Y|�D��H�����y��0�����x�o```��}/���T�V�$`��n�`��lH�m�ٺ^�D��q4�+�53��*�)�a~��)̒a�Yx�e�]����EKҥҝ�߿D�����E�,���ϿV5���)�1�5$�&mp��ֶ�Bv��Ή#�a�U�Ò��.+Fe4�`)��,�C�̻���l��iL;�x$H!bւ�U
��"�s���b10	��K�Ja�����_�K0��f�t�wLw�z���ʲ3,A��~�TV����[����	���������wmal;�ؑ�G2�(ᑑ�AEDDj .�� �����0u 2��F��k^���~�� �u,��i���(n�Rs����,	O#�|Dh�>-�_e�kN���T���p�~x?�yXs�)j<���A�$�욱���E�Wu��z"�6r~?f����^��>=2[5������l�{�P�,U:��������o)�iwW�nR�M��^�?{��r�װ�����Z�g�~���F�V�7���dy�d��X͉�G���D�F)�W�쥬+�~a��е�kD!�HՄo�BϞyl�}�V���X�S�D�9� z�y1̰���G���k�`"�A4�w�W�"K�������K�OP��p�9�._�U� �Jy��:Ɵ*_�҅�Ͷ��>��1Ln��\"�}�UDU�̛79�;^�c�4?q��q������_*��������V=�o�/+vE��D���aA�5m##�<.�+�_��:.e��0���n��<'�YKKk�L��>�70Psm��b�n,�"4�T��12�N�ji����=�b���xz�&N�\�wXQ�ųbO`�Ě9�<�#����2�O����Y����#%�*G��������~u�uV� ��>�|��TϘ�Pү��<4B�ߓh�����ڸ��EEE! �"5t��H� 7~�j����k���՗�@��8�뇊K�Z�}���[��d�WD��^����DلA�o���P��Л��S�*��-[���7�")�]Wss�{w�2^�rO��j+!]sZ$����B8\	:yͦ>i�AĔ+��^�<7?�DC��/<��`���?r�-h������s'��E�Ǐ�헕i���h
3˲���\(Ĭ�=|$�p)��@b�Ce�S�!{njzIS�Ta1�����0�ӣ*����'r�.��+�+y�>�E��*��c�ʒ(�$8��gS��!M����t�40����ٽ����&��[��ܵ#��''=��Z��w����k�7'��8���H���Ux�c�i�|��`�GCQ�4ƛI�(�n�_��>Jҧz�{�̜eל�@���swy�{���N�8�5�&�&CJ�Џ u:�8�Wb�t���PTrrv�mez�)?-�Bbw�r___�v�����y��C�_Ai��l�����*�Oi� mie����ߨ�űM0OЫ�1
1|dy�8 D�%�������y����v��bX�۷ʠ�?Dj&ƚ�5��a6�&E�d�uq���.4e��[O���Mi����D��2��:,?��}K��-w�����Պ�屎 ?����L=��A�01��X�<�%bl��n�з���ѓt����d��F�H�3�eS�v������T�F�ǩ����bra]�}�~h�`PO9A�zdG�qzl�q�b���n_-֥7�Ȓ������?�����Bat���;�	 o��('f�l)��i��49��?�폍��!������U~�;	�'^�����/_��'<�(�l��QTX�Z��v\���s��R���KZ����nz0Y]�Ȳ��Q����u����Y�q�q�"�ɲ?$�l��t$G�������d����Fc|�g�cf#Mj�>y�46�>���[�,�6��������ý�e�%�<e+�ˢz���'�h�.�B�g����+�����*D���:M�l0p�?<ݶ���2}�UJ�\xUoW���r�+��yU���z����]�B�86��-2a�5t��;M�Z��� �X!hvթ�IH�qA1<M_��,��!�`ǁ����!�ŉ�/]�[���j���3t�9�pL+TmG��NZ�SY ^�|]�U��
\q�Ɵ������B�t��]?OӅ�\�;��߫�6�S�����������h���#Ƨ��H����t�-�kV��e�����TV�]������.�� ��s�5��7���2d]@��e�^�W��ų�K藙���/���
�n��y[i�!u�X��׫���'����N���U�������g]]\�-h]=�SZJ�G�Zc��Hg:6���Kc;M��V�(k���֝�j;
�#z�ESN�~����o=�"_q+K�go�����n,BUEƠ*-��)z���$�Pzk1�U6�{,����k%�hoaq����j�"��#���;��e��ɓ��4�ۍMk���4�y�"k�R?DW��X��gW�����+��:�gYA��ݻqS3��8]Z򙱶v���f�R�#cj;Y�.��d�c!�{�V�H���f��BYz�<)��.譆�79�8)4t-�6�N��4�2r�O���O�<[SfX�OQ���CN�nߚ��Z�+H��&�w���0�":�$��LMMᾏ�+�⼢�:�d��̙����o9�a�L����W9ֈD��#=i+�I~�)�Å���[��*W�==�� ����L�S�����;n[	��L86�\��Ŗ?���zfm��Q�vDy�`��\^^ո������"W[$����̃y���˻�O�:��w�7Vu����ZY	�V�({�`����,��O|��B�G#C�3J
sձ u3�8�8�8���3?ފEn�ߜޘ��Xb���	���.f�K�Ӡ���3ϊ�;�M�{�l�eɴydn	�K]��f&z�J\0��S�=�}f/���s��S��t�� q�w��~��6�6��{��f�砋/����y~��rݹRE	@ ���D�����\�ފ��,--a҄F|/��}��{�K��M%/fƽ���A�}xY�K_�OA�+��db�-^1�g���7SXO���x�OT),=m���t��2�R�F�vq�kD&� `�9ֵ;>DI�!5�����?��ϟ?kQ����:G�ڴ\��g(��u�_��\��
1���o~�\����N?��Ar�}��p�Emde.�m���m�>�_� z�͂��*s�rN;��j(,Lnnt]s�jS�������?U��c^EX68\0(��`H���ٚkG��SQi�&��\2��~��$�{��S����B�aa*��|1�����ƍ�;��d}�$��ā������ki�zf8������itu$�<-M;ܒK��?��z`ˬC��QQQ��z/���ܷ�:*+9)�/HVWA���Ű�>Q+G�~�5��G�4 ^z	l�������u��F���M�@��y�...��On=IrxO�U�S�- �&,�I�:�mh����7���LJә�uc[ZZ���&奤� ��g�*Ȥ��9������^E�_�G�N�/o~{���Ąx�Ǐ!�[�S J�w��b|%�B�.�Cv�lb*�^f����Fg�H� D7T��]�]=�F_@Y�o��������a���*0�CSE��S-3�{Թ�=���R!��5���%��/�#%&�U� QW�f⵽/FYM�XL��:��5]7;ѻ	oR(uME���}GHC��+�z��M�2Ϡ�߹�c���qf��B����7��m�˗���Obc�����%�?U@BT�c�!)܈��4B���y�W	S���}�Drs����ګ���W�k�E��l��Уb���d�Ԑ_�۬��>e vQW�5Li%C�S/9���"�ima!<QL���_�Hgy���j�z���C����%XG2X ��yYl�w��G0J�:�#SȬ˯�c�ϟ�9�F���񘚾~���c#���:��,��X@$��2��4ߨ檫�#�����O^��0�;?wInt�
�G%������T���$��`��/_:-���]jOI�/�wOyI�o��Ϸb��@|�ր� L$�v�J[C�����q�����ot��$q�1���UH0s�$���Y)�X��yӂ4J�E[ۉ���{��� Rl��r�͓�"�iߊg8R���G�u=�aaa�/|���D��i�"�ɭDn�z�)+��,���^��L�s�d`Ǖ��ﯺC��FF qpu��շo��-Mj,�b��5��jmu]u���&ǰQGI)��]*��� ��Yj���XN��Vv�g��5,���k�Dq�T�V1����Μ:u����(QO����Iw�h�e��b�|M�������Y����u�f���U�����9=�WNi��pqs+v ���ΉC�|oet}P����0;8�ƓL��/���kp	Hj]�f}��u��������&!; ��, P9儒R�8w�]�CE?�+���ʊmv���=:_ޅ�B�����}R`�UgyYb�d*;��|�-���t��k��o؀����8��p�;�z}9+0/*�g��8���NW#�Ci����{X|���m�7D�V���}p��{���	��������Ĵ�J��������{��ڽdw�r���:+E���5=��p�:	)�"��	�����>XM.'������{�.`b��J`l�hg��E,�{	�����KF��;�K���������1��Ȫ^��BÆ�@ŬD0�0#P��G��r�_0G��^�e�\i͇�x����՗�(����֮X����rNy˚�AAA�	�G��3gB8v�`g=\��\���� ����,�]o^��0\8"_fI���W
k��͒�����qx��-�ϲ�-�ܘ�!����7P��`-��tg���_��X#��  ��fxɍ9�[�����Ż�ş�G#�>|؀]L�*��?.=R��<�+1�6�����[&�1Օ]%?��V�jݶ��K[ �O�o�E`k��lc��2��;*����x4!��l�������l#�n�cOpGd5���K]����V	P}��y%��Λf��5�v���#�����`�߉�>5X~��H�|Q�AB���}`��'9L��0����e���ف�$?{���A}������U����ϟkCd���{��@�
�;�wU�<��]��~���A&ң�htWOX�D�ǘY�3���������h0kj��x���F��|ձz���Ps�ҍek`�]��x�$y�Y�ğG��_w�YJ��v`�m���z 0�:������}q���\���$��qC9�ƏO]���:?��{��Z�u�6{\1O>��W��4������;7Q��Ӑ��u���Ȫ@��{���V�L����}�ӈ^��^�0����F��%���I��%e�u��#��2�Y|ꋳ��O�N������	´�����J�9:����!�����'���F��6v�eK��^V���*�]p�&&1A����c�W�S6�I��-�%.D�{8<))�g���r����e�xpt��}���"������P�)
���QX������y�\ͻ�B���wK��yR�u��J�W݂��w�##E��{���Nz��Fd�?{��Tߓv|x��9m]]<r�I�'z��u��
ּ�h�[���8�}���X9�<n�^�﹖��x�Ʈ��� q�� ▛��OKh{�V�C�B�/��������_�l+�Ni�4��Vd���j%��C�1�uʀD�i��{Ί7q����~���C`��[�����!pb5޺�'NL�,a�P�L�����e�uFn��B�8�2ȇM�+�Q�nv���d�-�R,��
-TnG�@�����c���w�<= �(��{a+�i�M���B	ݬu���'�G�o�|xZ����r�5EZFFE/RS�[\V8mCX�nɲ�X<Y3}ʝ�-s�wuqq2�t=1��RP(
��r(Mxaws��ꛚ�A�R*�v�`-x՟���[���6:{Z��>������V]}����e�,�[G�WeA�����&�ܹs/ �����a����U<;o��L��>MNV��|�l�vc�C�C��q{2��{ݼ��B.=]MP����gW��ܺu+���RpU�������	Bܼ��9 ~z�0yuos@_�Ij0*ts>B,��zx�.`��& ����l�f?����9c���Ny�V��8�Y�&Do����_B���>�;ΜY��G1�?&�Ǐ� �#���6�FX&�FP���+��	��|+� n�$����6�.	H�Uw���/n��]�w&���?�F�K�t��ؓX��I
oa���z��9�ѭ��7.�T��S^�,�NG[�A�ǉ1�8�433��4�|�dxu��U?�2��*C��Lyf&O#6����v\h��
��
H��@�SӔs9J����(�8=R4���9m�4{۩�z�їͣ�]7q�)>�XOKU5�J�ψ�P\̦���C��S)II����t�;'��zY��fQ��֟^]����%O3vC$����I��"V������Z ����u�Kl��C��i��W�E�nɶ
�Ld��o7Ƴ�\�@_��;9+K�'�U�P� ����x	� n
�)��F]%%��m��
d��GYQ幯�%� �X}dU�����Rh����2_
,?�XҩѬ(�����m�]�.v��{t���=֑�mm����/���QL6��̃X���q�"P�I��x"�է�ֳ^s$h�4)����5��N��<��R�9�K�-Ln�m��u� 5ʢ�v8��N ��o��{�@avt�T�����h�c�����A�.q9�s�Δ���� ���Rd�Ӣ@<���].7���>T��6�	H�?�o�c�Z�5?f'\����XC�Y;)����q<ڕ.���f6̟J��n�LHY�.^�+z.��w� )-�@4���̂_}]]_�}M[�d�k�
�D��df�͛7kkjnU�I�sS:gcm}�dq�s)�[
��	���l�V KD�^.TB��\����eom�d��́onv,���R���O �� ��,f+��OJ�}H$̠6�]J`���o�����	8L#�¬I`yjR��t�O6��.Yn���RU�ޞ
ԃ���0�1��z�+ڶ�X�0P��յa�C�֘c�`O<�fkm]�����ǉko���<9���Qgz��� d>9�@Pd������A�v��d���#���.��x̐c��m/M&�:��e�8_SWЋ�����Y);1�s5�ݤ�/^��9҈P�+�fz�74���ٽ���*x��Y�?ut�(|j��tކm�C� K�zr�L2�b����hƖ8�`��ٮ����uo��Y��Q���T�7���C����G�Jԡ=	�n7ဓ�`�����Ń�n�	~:vyzR��~��ӆ��c���N��66����"�6�.�R�'x�E�}��D�4 ��|m���C����/�h����57��Y�j����R���&D�Oz	PYag�WL��*�,������i�"��Q�l]� O
���h%�g�e�]dS;:�E����-B����9d�7��n�9�ќ��v�L����@1������6e�s�oq~����5�X h@�0���ଜ�|�������>���P��x�)R�����p5j�T!:wUa�иһ�1�|��L��� B���a�!H���a�]�o���:��U �2쓓�ٛ�6�Ra�0�VmӶ�O=����-�I�d�<>}2''')55��D�&v�b/�R�{
��/��/�B0,p�8�H���XJ�F��:!�h���}v�W}�љ���pC�o;ck�A��S��۟���v��T�;�.ΞL�%�f�މ(�a�ܾ}����K��M���RX"%f�G���P5�����/]s[�Q�U
l��� ��^4��t	D5�y�Й	:T0nɂ��EǮ(*NMM��:�ڜ;'�j�U�#�{�} �	+e�u��"F�8�f'I�.�7o��	��,�,��
N����筬z���{[�4ͱsѵ�65L��55��%L1 �=W�;��?`oV�b�)""�K '�͘g��+LM���{n�D�a�#�6� �hvvvxMR����4l,Z��}8���tG���W����)�o�����ʒ�w���eE�����l�z�zVB耚��P��]���du�3��?^>ć,�$�)r�l��������s���G��NNHP�<�!�F/"ǧ"Bt����[��6_%c`�t�˅*�{�>lX��$+訃�ML�qe�Ç���S!{���5�;���
(�E�VXFw�i�{x8���!�!�3��k����P`�|��F��O0�h>�4 E�/<����P{�۝C߾�T���6:)U� ��F��9 �U@�����,�!����$�K�lCC0�˽�:�ֻ����Ģ"#��~�/bt6E��Y��Ƿ"���-��冷!&rh�$п��B���\�
��Q &�wN�da�EX������dߙ�!�2����h߃��� �jb��G���U'��T�ܬ�y�f`l؂J_�A���2A�v?(��������_�<ɧ�D�{��|������˵rV�����(sz��o�(�0m�-��bߤ�t�Lnj�x�k��r��<����Խ�FY�?�����k��#�AE�**D�F4"D%�(C�B�J�$��d���E��!�v)Ҏ����V������\���sux>ϳֽ�{=k����گ*�0�(�����H�Q�-p{2T�p���er[�	��XZn��'�$YXX�O�I��;3d�a�l{��)k� 9��F:�F���r���8� v����`��%�_���tl.>7�ZQ��Bv{��D�;��*k��nG�bmI�W�3=��8�l�B2�!Gl��d�YRc�h���t �K��2��_mb~���NG.e"�rrW� �+��̨+� �������՘g�Y���k ��'���ssrХg^|W���L��(+:��^ȃf��6���m�V�,6@0�b>����/�����LMM��aK�3�q'/����N�� ��f�m8�����}������GW�{��E��fi
�1ꭆ�k+���.������Z��%����<{���'�g�C�<0�ׁf�������o;>���?/�FA.�?._���U����+����˗`�#LbC �,���)�m�K��L�X���ÂƼ�b������PK�fs}\Ⓛ���ӊ�rm�V�m�,[��
��0��]'%�l|qٜ;Z-���msj��#T�f����c��֌�w��YW�Y=�ۓXPp~�ݞ_�w����M�Џ?BRv ��]���14�h�ڻi%�bQ��+�}�f��\�r��0����Dh�X>^$���c�#�Ve��͏��Q�MIi��%��n� g��7] R��Àق���(���:OO͞�e"�l��D�hg���q��6?\*��wH۷��fs��=�us_�=ۥ��L[恱m�`,����G��rY.3.#������u��)�~RXh�%�9�ıQW=����^��)P��Ç;B�4��26HI�򜭍��v����_'ىΣ�v[��6��[t���X��[�y��X�����ْ�K�Y�'U�\zJ���v�����~�5�;�J�ir��W�lr0���Z�C�������PP�D���m_|��$���o9ſ�c�dz�	��b|���������l�t�������(�"�! VO4j� �9�����9�~�/ׄ�
�\������n�����-g� ��l_���Җ
�ZEPK�k�u�M�:9��2H�5�"Q��S�b��ÜhG�ď�t�Lu�-TJR�����8�ՠ�����0���ظM��������J=�k�A}��
�]ۥ��^�U^0��_���O�C���eNO���s��*�ǒ��?�����x#J��<�0?��\��2~� DuO�M̀
.�fϵ)g�X��	���UUU�O�>%VXbf�wzw�?c��b���� �`��y'~R�׏��V���P�>�C�?�\R��*�Tl�u���y�l��ŷT�l�p~�A{��EDD���a�,�h��
�k�i}a�6l�j�ef��ߪI_�N_-,̨��wa�Y�/�~�'���k�'��$��1���R�b�[Q�>㈩Q�s;+~M�Q%�C��gk��y�ȋ�̃p���@њ��`߷g;���[�la�9نhY@f`T�����/A�
x��ث���8*��%p����S�3v����]<-'�q+��4+�We�ް �����+Usl�yKKq�^�{ �T�7���: ��Q�����U�qn}�������i��ȸ#e�㮩�g;8Q�C�n����� �f���W��r��Wճ�8�-:,��s��a f9�8~ ���.�#�Q+�7����fmڢ���0?88�o솈��`$UwT�L�����e��"���
Zon�_C.* ����Y���@�C����æ�rNNN��0�	mXG��@C�iWܰ����9S" �<�>�d=�`@�8��?1ˉ.y(
۶=��>/������yم��qbب��*���ҝXe,�~W���nȕ>�՘}�8L/�� �Rlj�d��B,��[yZHJ�K�v��u��YZ����|���OW�.���^(�ԝZ˩�.���~����P����vc0�L!�T�.[�T\l�s�<�4���nj�xac|X'�+��b�,�p�~�>]���F����2/����*C�gT�Ӽ<x0N��+#����1{� '���a�A]meı�bb;�#�U��������-V,��r�Á���%d�Q^^��>�eUM��*hN@�n�_ꛏfP�0:�ɭ�5����ߐ�:'�������FG�c��5;�W���pK �N?��Eqڡ���^�"IK9��ZL'`n9����ep���˰� v�ÿ�3���{�-곗1D�"|������>��V%���� ����do��eW�"��u�7px�k��A��>�O�w�e��K�@�z�9r4���k��K�"��]��  �kbR�e�Guu���]�H�v/�"(�|KX�G�|�(�~+:S�F��2�����Ox���X���Z�QK]l�Mojl,ߠ�7G����^�:�$ʀi�
Ǐ�^}�ںA���K]]��v0:���~�Ui�9��Q��LԬO�;zz�?	����Kj}Eg��!��c�	�]��\�>�:'j� �_�8�]�f�)_~K�Q�$���jŹ#��A��=���#_׳Ҵֈ��l�j��d<��\
_��R,�D�У��t$��_�fp��ee�Lvu�<���]�ҩ�X-(��W0G Q8�/���ġy�(р;p�^�o����������'�[��!���
���(f��n�i_��oo�&�����[��eÕ�����ȡs�Zl���5�o`����=����	�Hi�Kg�/tj�5ٰ0P�y�F��M�5�e&���Z�X�"��۠�Z�TjZem��xo�h�xl3>>��ѷۻw��8T�D���c�S��)DwP &^^;~�������!Gچ�L��SS GsN5���jb&sw:0i�����I�u��l#�����'����k�g�+S�����V���m;v`�{=�h7����A�b�o�fO>���&|��C7�3�rą�4�1Y�Ծ(����=����?�
�!a�t
doJ���[r
d�M����W:n���|���Y�ھqY]�ӧ�=�(�o�Qm�P�?�����ܫO>���
C[e�y����g�=.TIA�8i�5���nm
@t��ߌ��S��K��g
��Ҏ	������({��젃Y�o�w�r3,l�=������ߥ����l*7W�nLF8pkӍ�{����În�=�vM�+K_��{8�0��X�pѮ�.��^T���Dv�>��M�gδ���!�h��_��1���`)/¬F�2s]�5�$Q]� PM4߾[~7���S�Y�#G�Il5� ��[G���4c����OH� Μ�����-�Ǫi�x����_c�p����K���(pÁ��">�
�TVW�Z�d�dɯ���IFv��.h�*OL�b�g���ߋ5�l��|��ѷ�-1�V57GtC`�3�Q����S�&����J9+����:311q�`Wl)콉�C"���� #pr���-��!]����`TsT�%Tv/;�؆IS�f[�����pi�ǭ3[*��@���v}��O��Ƅv|2U���4.����Wr�t���ׯ]\Z�xl�4��a7O��9�-��߿��߮�+*!q�C�u���Eۜ�����Ě����e!Vƥ�mYܦ��ٰ�	�O��n?�>��������[dp*~���C�AE7�����#O[
h��ن��2W �&�Cm�W��ը;�k����u�����fF�m�X����`m���t��$��yA�\~���֭O��q������%\^��k��ս2228>�����W�tt$/]�E�{H��9���U���Y�g��.şs�=�@f�L!�l��F�8`x �q��f"6�q��ˮ������)�ũ�ʲ�o����UjA��:ur�1�J�Y�,�.a�ǰ�8Dm���s,���I�)���H6�b��W�*�:���uj�a�f��qH�����IX�[f��Va�L�5@��'O�2���� 8c�^�K� �F ������J��j��UQ9M�\���}��?9�Q�}J[Ugw�rq�%��v�B��O�0��w|е�f��տ�~]��I��.��C��ž}��bw���4��6���L�5q��-�^=@��|j�P�sPpM��3��0s��ƖU�%�H�~����u.3y�uKX������'$UՖ���ǪU���q!"�9'�y���h�ZZZ9Nm[�G*��X�[U[�rW�� oꞰ��4E�����uLR�,������9?u��Q�㕩))�������ViM}NV�
'��߿_Й��3hM�)_w�*`-�(�KLY��"�7��<��#�>�b�'�***ZU����~/�G�@�����qqef���n���"++ٽ�����`h��_Ɖm�R|��,�-�_�j��⁊G��]g	/Ee��s3��.�5�����ws�vu5���Mh.p��Tt�?�kW ���l���F��,�ϻ�}���_�� gU��?�ᡢ��:�DgzG�|!y	?x����A��
=���%e�S��?����GDDĻ)�|�j')97�k#����������X���������8���-�!(QGLMc/��� N�=�!2�X*�&������S�jH�
C����܏���
0Р�u��%�t(� d|���"�]X��!�@��rU���S���/��/���򪲦�����sSzzK+\A������;�����Ç�y	))é�5 �AT�w��1)))�q����z�Z��I�R 2�r�����C�*���(�3�y)|��z���I��߻�?�N&½�ܕyk(����{�o�7Mب;?���s�@������;Vr~��!�)�a���kuԜݪ#:�N�ݏ?�@�+�K��Ӽ�1������	án���KJJj5;�c�M�1{pOκu1�j�F��G�D��ɩ&D�R�M���r�4`/5�������w�Z��*w�� *Wm/:���0ؑ߀���勭�h��V!¶�y��XZ�l�]��6n�UU��U����bp*��M�54�����&à(1'G	�龺�'~NO��]b���%P�+Ae��	z�S�M�ViJzaZ�ŋ����pߨе͠s�=;���X������/NC=|�.$6��V��W�v�w���$�10�9�}}L,��`����{�y"quS����d��M)���+�V�`�F	��Swwf�SxY�����'?~�	����6����F^H@>w��f¦I`����Y9���E3����!r-%;����:ߵ�r�Zuuܰ�t"�E>	�0�����o[�/��A��[K�D�733��x��gK�����bS#h�o��TѥP��Ć�3u$�+���.�z��p���k��wo�~g��	h#�A�I�{�	����!1�C��\j7>$&�����ֶJS#�t���K+'�E+��"qNiCXtCQo#�`G����"�N^� �Q&z��  j��vo�A�V��gedI�ۂ�ץ+ؽ��{���p�sA��п��V�(ې��ϟ�|��DߗM��x������x�X��<����Z��Y�!	99|�w��n�S�����zzo?^����{��f��**fe޹*[��7:ӵ~��ϯ��_�O��J�b��;��,,R@�W�u�Z�VL����X!�f�r���>�	�j���C|��1x�ki�:>�I��ڍ�]@-�gfȳS���pO�i�"���'�٢�=�m��7�����HlQ|���'XU���~bV8ic��Q&\Ra?jk���V��+"�GG��ؼ�@�tk��d�¤��ә�kx?� y����'��{,x�5~��;�Bb���|߿H�I"�oI)�y%y�5^PP��ޘ�$1�~
��Ĥ Wc����f�D靻w�������Y|~�Чj�O�W4Sf*4f���g�F.��õ�ߌ�hf�5Î|WS�;��K��-/�y�&ˀ� ���Cc�iϹ(O�U�7= Z� ��|}���nӋ���MVvv��mx�2FM��GINmiX����]�1���u���E��&x�0:z�����D�-^��߃`��MMOO)9F��G%$l@L����m�6�����*��n|q89"22+�b�ͤ�
��[Z�%�'�*nz1$R�Eǚ4�yv͞pټ��5��|_q�}%�̹_ݩ��:��AT֦��VK6�����1N��ӧ7�U	Mp�O����0�����T�H�jB�lkoOZ�d���{�����w�w�� �x,�A�ZF�ګ�wc~��B��ye@+�T�g]?�?R�I1��=�{>�Bt�}���*�3���0Mb�#[��cM"w��ӈ��8v�8v�X��2��EF��� ���� ݿ-R���������|�'��b0�DЖ�W�� @op���/�%2mݺuH��Ah�D{�\΋2tb~��/k����;��0v�~YHu��%�G�ɩ���[����<��yi�8��ݫo�'��xVޟ�,�؜u�t����!���\�!�{޳���'q�ʏ����c�&DϰHØ�ѓ�Z66TGUQq1�@�����&�8��/٨�B����U=�������.�Ȇ+�O0�FT�'�F��~S_�g�{v��x��6�z���bS��V]����vg-�Hl�ߊҮ߸q�JS�&�E-�������Z:|+Z����� ���B
��A@7�s���?�������'��15�@}�`W0�\bVVb�A���ũ�2
�6��}�O���Rf+X�06�9X,k�:;;�S���d�R��1vu����_�.�>?Ջ�d.�4����;j����;0e ���$��\dO2�7�ڢ�!���و�7\��ȈH`�j0�m۷�5���
	���N�������Ѥ2���Ý_��U��{X���W���ԌÇ*�y���Y-"�k�L�md|�����b#_<�.`Ӊ�N�fn��o�m�����_���c�����/W���s��wG5����yy��Ũw��(�ĺ;$K��W��p}9�U���{]]�����7o~7-����Ξb2LI0�M�'�������97M�r��&*����IYYM`ȩ޼�a�>��Zq�֜�)�J���M����K\�EK�*�/3��V��"�5|���p� {Y'�u�f����/�0��0�����Ni�7�`������	=��Hgٲe/������bMB|/2M4�D�ek��Zd|���%�FF:�?	�岦��)��T��u�|L����,q�|M*� �d��-�d2�������!X�<k�O5cQ��;�>h�xQ"�}>B�+�;l<�h�����J�38J�i�w]�v�fnn�Sy.�e�}���v��b�������/�`O���2NW\Y�`��2�����m�T���"y����=���մ�I_�(�]�ǼR��Ų�r������~CL�U���D�md��3�z�k�ʥ�/�|C+.`�F0��}�zUAZ2Vᵴ(	H�ҙ�z��G���$7�Ɯ�����g��M��`�\A���E56���q9Փ��˲�*���hK���U9���Tm"+l�p�p��!SS�y�t$^�LLL�a:�_+��W��[&; !��;��Kp��~�
�p�b��uuMGn~&�*��f�R��V�(	�������"uq*;[��g�~������[��� r�l?�U�j����>��*�ۂ�==�@_ ���|��8-NxuSU��Fv�c'�V��z0|Il,�BF�������3��"$ϫ�n=Qŝz4�ⓧ�;��=1���q�+�+�c�_�?f�L���D�r�����;�\��@� bU������l� ���c�*$�ǲ�B��D|�������`��[=�f��:~�$��L�I}��ï�����x��w0��h���&n�``㠆�9�<�G�N5�S��x��~ae؏��Z�T��+��uAB�u<P��w� @m��LU^N~N�F�L7fc��-��M_ jc"*Ћ�8UuaDc>� �t����^�Fn>��GQp�̟"]j8G�e�q�YS���ad����܎�Y'e��3�<������>�1߾�읎NH/v�::;�PJ��PF��6	���C�G�8=�j��d����훴��6��&�$*�H�їuq���
v�H6urJF�.<4tx��X߻l�퍧<��/�%����Z�^���F�\]��3LC�qq{f&��SMutu�՞tvZ����b��^B_�����t��}(�j޾�Il���)&a�8W��w2dY����g����m4�i����ԟ&Rx5���*U[%22ޓX(�A��/�Z�땑�؊�5�}�y89�H�5fx�X�*�ت��k�n5Hr�D*0�	0L:^��_��K��Zo�������l�ŋ��.��w��?���7�y�0�������Y³#H|d=���ڳ�A�#GM��p�^4=�V�f#��ɢ5�pԚb�Y��nnñzӥ�0��<}�d�3=I���~8�M;D8����\	� ����'O��ώT;g���
b�1b`ԡr#삕�	�u�c���LBO���ի���u�G���J�������X����(D/	�ʦj� g� �Z��j�S��E��Ƈ��S���e}_��-�> ���.謇�#���a�u�TL�:$�<� �7��8���& ��	|\����Ŕ7P9 ��� a9"#�e�(^����kš�f:z�2���Ϥ��E)�),,$y��$����H�%�0�Bփ��4L���K�Hyꤗ�.�pMݳ����<����z)�U@�O��n�����9��}��ҽ��Y����655��j�����t��}0�c� 
~�P�"t�{c��v��?���Mn#��mm��R��Ilw�¢����ŰdӣE�ȼ��L�m�����Z2���}o`f�﷉6뀪15�X�飠�E}*�2���hk����FF�����hM���(����$^3��U��S�@ށ��2�a�DG�0��X���s$A��67z�a}o�%^S�sp�ޑ/���( ��J{2��hʬS��A�-�E��c͂��)�B�'\SX(�*~Sa[9@D�Ȯ��'��q7�k�R)�x·��X,�'^?����l$��[��U�����s��6@��-�͕U��2:6v���d��!\2�"����@8�]���)�+����S-
�%��3���y�3y4b����Vj�E�K�Sk�WN���߷L4��gz�5 �$� ���>R�+��D���F3�<z$��,**�$6�>�՘G�'z�����Z���m��k���1�~ǿ��8�D�gZ�L���9�Z����LTml�&K'KxSU�?a<�����%��/��91�Dx߹��ǖy��) ^��,>��@ǲ �0�k�����:}�@����;%�;�(L��ܦ�ֱ�&&h�:޵��/���ʚ☌e��G��_��{<Nl`z���jm��&o""�W_;�4�*����K-����=-�ʦV_�E�Q�����1�dC���F�����x����6j�S$v�ڄM>�Oâ�0cf�~�k|�I�d�}4��C�(���pu�X	2��m���!��ˮ���Qߵ5�>�-7 t�b�w		!r��xu�8$�Ymy�,�ԤY��T����j场ۅt��9��i�q@ �E�'^�OsqImM�|K��o`���kArL�(^q���{a:	�=�Yű�_��@B����������#�?I�#��hl�<`�+ ��*9�UAVi��G)Kh�6��/�e�p������@љ޻�w6��<3Ԙk&��z6��3}V��fǙ��q:��zP~(����=~K�+d���n
)���/]���,`�c���ȕ�t�M���tqٌ*�7ޒ���ޝg	

��wW<��1oA)1�׭4���W�k�9mZ���5�>/;��"6�:8�����֕�$`����TP
�4Y��M��9	����\��G��Z>(7�X�l&N��r%�!����s`,#�+��#��Oz}cU2�A)��P���K�~�Kzf�K&�}q�6��K��e�MB$����Rn3� 1gB_^�2A��z�k�M� 8�8��F�������Vˋ�2[��캨?�*�HX��9`�Wq�B��:���dr.|W���O���v,��$ԉ��Ʌ�����|�<�En�[��|xq�����P��qB��)&��5�""�sb���@
8�ܭ��}L@l?m|4�>:��.V#l5	��[[@h�ϴI��<?)��=�?��k�������H�����֏9K���Uq����S�PԘ����T�>p����~�Ϸ�:�R;;�H6M?"_�.��v�z�'G���?��: ˲M]R���m�)���7�XY�O<�ݯ"�԰uu4�I�_-���hU`��(h!6b�n��:Q��'za����a䕄�3 �`P�|��¡0�$�u�7
[V���1sd9#Ȋ`I2�qf=a���3�1��z���{W��%��a����r*��p�谆�US �ü��!�W��>R-�*����,�YF�տ�'t��G?Ƨ�Y��A����� %^8i�.�&���xayg��X^D������x#F�����¼|�Ib��F��O�8�&S��V���O��1=����8���׎���;}��*�$
�V��$|���Q}�	4c�u(�����;Α�5��1���;�2�fj{������Vw!A3���l��~��=��Ǯ�W�{ݼ��J��F[$YÅAKWmfR��E����� +�x�<�3��r�Gl��@�b��^�IG����e8_��o��������}������}�T�Q�x�.�U�$����'2��*׋�L���8�U{+��9�lJ�"�N=���S#��BaJ�H�x���������8'��Fl�ի���q�Y-�hc���HL+Hl��W`%II�m��������A����X�������D���k.����H�=�_�~��M��p��>ji+�p�j)N��~RZ����y�A�l�>�U�w+��s�۷�5,��ئ�d��_O��IV�xX����yH�.r��mY|�ֲ�XU�z'��	�s�"�a\=3�l��EI����U�>[��H���Wr�|�������T�?��;t�`K]�N�u��C� ]01����)F*n��i�����2J���'��] ��3��W;�&+�`�8�djj�	�O^��S��@��o���%��z�C���?O�7 �~�`�Ya�w��1�va�s�7pRX������tGS�i�)�^��t��)�U�=�EX�rN���a�]0C�H��z�&��9�2�shv�Y�O�����z��et�la�S�E���:?��� h �*�[,�Z��;!����^�W�������@N��m;���,�^TI�J��o�*��S]%d̡u5ZX�<8���K��'J�@����ZR��a�EQ��xD+�OHp����q]��t�PW1�ٜ��!3$7���%&j���/V���o߾%��`X�+e�D�a[�CDt�����.�8A-��E]��4��ş �	��CulsE��a�p"=���Wi��Bg�0�S��: (�DX�G�] �d����Me7Kq	8��$+�cXl�7�Y�A�����}�d3�c/����C5�?2v���+��A��aD����6�|凓�-�V�V9{�a�ΰ���Vӹm:���27�-MoKw(Q�TW�brl�/P��7\�1�Q6g������C�>OJ�%�Z��V�+y�鷴�y3�>�����p2���.X�	B���1&��B�f�S��f��b��n�?&/u+�*��FO�u���"�~��'%tw�HN�K��w�F�����X'����82���Fap��D�)���ٸ���8��Aev����Һ@���Ş����V,��D��?���C�<���y)�HӉ�ᩪ9�ٯW�̘��WeH,�AAAH��0�=,Mqؾ�O!�K~ˇ�&{�\���U9��#��g�����Ǐ�6\������+� �f�6¢>_�K�*��藖�nK�;�K\G�ӗL�֛��΋��� -��Çq{�y�$��ȹ�-2���Ox%����X����'03RT��6�?���ZZZ���@ ��@�����֐�],l_U�}RP~�����c}ؘ�@�K$�~��x����"�yPA~����ӵ-!���彆,0+
�f�����$JA�����E�J�EB�Jt�hz��I,V��l��ŋ��ٯ���*=��6z(�Qb����������I��ʹ��n����҃$�ۊX����'G���F��� ����y�P
���b�ttt����~	����3��%U��}�1)B����7_KKm�r�M9{G����>�cB�X@'��,��RA�Q��'n��������B$�yL������]'���$��̑㩨�a��G�]X 1dG*��!`凍� `����-���Ӏ>�YS8�s���.C�y����^��M��~���l�wsVm�ox{�H�޸ƅ�"���ii[B�G!jz�s ����AU��Ϥ''g0�,_��:Ɲ`����pI�5�{B��Է�X��ۂwDxQqqKS�m4�͏�����oܷ�����m!���k<���:�	��PE
�G����~���90�a���X��y�^��b&*_���$�
sߩ��5�ؼ2��!��D�.������k��_�Y��̗ST��c&��Y���7Ě"[�z��q��:�ڣX����{6}�{[� 5���r�ݔT	��xc�����T�W�3�t>����~��f��vI�����@&�&7���<N	��l�WY�!7,��?S�b���s4�~A|���#G�t܄�5���l ?����`t��m���6���������g\<�w����{��4P/��wm۱o��EIN�𖽲�E쌟��5���l����m���UB��v����@u��H���H��#�� �>�_�����~ꐲp+�W��n���۹�lzjj.���g,����������E��a��Y�1:�\L������2��W�X�����14��N5��|��ܼG������ƍ��G�A��tV�-S-����.nh�h��nU`D�W�sW��]��4�����w�p��'�m���%"�Ǉ:|���-���.��:�nL̙hf1o ��uKށ���?~��As�y�ѣ �/�>�x�%�΅�1�%(��}b�vCk��[g�B(�1�
ڬ|7��.�"���ĠTS?�q;�.?��{N�0����d�����aV���T�����2!��6����PG���������e�c�"���+Wp�'#�+`��kV�J�H3�<h�W�/�Soڳڻ����5ׁ��2 �0��w�hb�ai�W����4�Ʊ"�$�y �e%��{�n��.a+�y:�^�Orz� Dd�Ĉ������h���k!���@���Y��c�R�t�$?�QO$p�qb��c[��<�uzJk�@�K�1%�za=t�)�!bx������T��+7y��o�0	�S
|�������
��kqC��;�T��4�"��?��FDDl�d&K����Z�J&y�\�s�����ee�R�*�q�3��t��[ Ә��;�� �+jG����C���.�G��Ƞ���w�v����
W'�z�|�hɨ��2���ZFg����p�͛�tV�7�L�Z�#G�cbL�і!�Yi���$��c��Q�x1	U�RG�6����r#�}���6�����!E{��˸���Yw�G��M8X����򾋘v�un��eЖf�]O���Ƹ_�:�o�>��(#�9���3�ĺ
~y�a�苂ٞ�p�W}8 �C�W�p�x��I]o]]�O�Yb�7�D1�(Dl����-�I�R��<���]�/VzE<�_ZNN��l���������ǖ{7e�h��99����vq3.	J��ʄ7�(��x�q��21��zzzv��9����}��"F)e4�������W�_�)b)��{��RGb�7��:M���X���!,��� 6����TBND_��Ժ	d�~M}lK�Q�Eʠ�s{�[��RL�VOLDF~���m/Ub�/6����4ɪ���R��K�&�
t�����<yv�`��S�ΜI����C��ف�m�JD��ۀ���_�4�-a��8%��iO�f�+羸���E��.���6ן>������&x)Ⱦ���њ�H�S@�y|^ܹs"�"+��+8��.\����D�l MQ�-JR�a���a$W6�5�E����
���K"E�^���X^���������әT���L������Xįh_�a���8�ąq�xU�֭[��Iy,��<�����a�I��<��g�]/SSc㓿G����m�0}���4�����k]�4�*���"��mj'ᶰ�)YX8��>=}�q�*�s v��+|��|v;���X����I|�"9Ap�^��+:7� �Q��Ow�Η{��� �A6����"=&E�����Dݳ�L���������@b�-��|)�/�W�B�8A1�aQ���VN����Z���e��55W�!�������P�?�z1�[N2��Cb?c����$3Si�!�<+�/Dbㄅ��X%�u��Ԧg/y	^'� L�M�?io�h�Аo����D��=^q�ƭ�=�� �W�Z��"x����?�t1u�={���d-�?�Ig��(�QCvVTD�sK<oj2���na%��;���Y|H�*�7q���@
B"�6�/�ʚ�XL��k��}�$D�J�W���s���5��4�s�0�B�D�(m���gK��Kň�7����'�t�XZF��w|:ǎ=`dq ,�cJa���@~�0�9/�ƙax��N������lr	6`���5H�a��"��l�*����JHI�2h�p��M�#)��̘NEL>��̴���S���EOd�����}7V&�f�||�?���������ҋ�>�e�����
|��<�1v�w�S���+�N�&>KN�18��QFL���"������������%��Am�>�/�~�s�藍��{�H�mdv?���8�k�Z+(��#(�=z����� (V�=+�?��^����!w�9�·X��!TL�Q�P�/�{)��͘�DJRrD�����eգ�	��@zr\{v2��_X0~�����-���� ر�<$���/C���[���ן��>�iz����
:w�s����4U���$�����z|:.�"&GF�G3�Lw�f6��.jյ�(�4��3F��B(Ђ��qG	t�>���s��a\���wc�B�_m���*!�-EL�zz7��C�8R�)�xh���.3v1*�u���2���VIL�#��YM��p^��fO���}���IA&B~�-�\��-�ï��0�7lw��r8u�V��d�	,|y��~�E��ËE�"vvv� �����G-��髷�x�W�ii �9�#�7j�l�!D�89%o�.eTU<~�H�ߠ)K������[uK�as�륏	#�zU:����������5Zn��Nɦt��|��K���:�M����G0Ҡ���ב��!��'�b�N=]�*��>|�����bсx�OL"�D�5��߈�u�woܴ�'�p����`�P���O ���S#���$���a9Z�]��v��
��Pݚj~G�a�5�)՜��jF�U`�Fi��	�n�L�,�BT�t�vjKk���r�V��c�^ m�^N3�okm�ҫ#�ðį����߅�d��=KL���+����i�-�m���P�|�(�������rF�5�y����cU	��l���當n=[��!�~J��ĉ^U����)��KS^qK+���P(���ș���,�3�T?��"��7��,	ڍY�8(��_P��" J1܌��@ N�Yl*"$��:;S�<YK0��M���K���R��U�c/�ԖS|g?ي�g��,��OR�	�q�} *.�]QSWwDsVVV�	e&(i�1%�s��>F�0B��Ȩ"
��O8b�/�g����L����Mi����
��6��U1yyy�/X���VwM,����ѽ��<��G�/�|ŎO�>��Rt��f�����(7�����q��ʘ���E޽�3FT�ٝ� .|���������[�ސ�S���f3�ГLN��m!�h�ry���'��w��'m����ʈ�"Q�ת�RY(�������.�*Ò&�K�5m�����x�
��Gj|�:�V5y�"������U7�pT�ٳY����= p�cc�2��ڡ������U����ϭ*�z}yYnϖշ�^��~Q�����%l�R�?&Yb1���;/.�;���D�d��jR�Lj^�y�I6��S��v��#o�~r�
;���u��
�\
�>�������_}Rq����y�&7>��V����t^Wv~�ǽ+��������')����������٫��zn=�"��I���`j�V���I�ZR��\
tARR�`$>�1^! p���������m��Z�����{]�+�.��4�;�<��N,�|E�O�C��f�eqv�w��X��}簑���T��&a����3��I��W(����`�$�4�R����*v/�Ҡ�kQY2�v=�be�	X��,�u�D��`G��ǈ��\0��	����\�r�Blǋ�\I����V6�"�� �� 瑲��bk
.iL;,��U��k{g�j�ο�?K�ќ�2?/e�(���,O���VjH�s��
`�@�$���!0*����J��16={�L����aq�ӣ��]�q�U8�
�o�~0��z��R�W����j�q�z�s&qf����x#�^XnIK�g�L�qh---�BWM��۱τQ�&@����濉߿����{�elKW>G"��V2���a��o��?��*I,a>1��EL��p^�@h��K�t��
���Z�!4Y�>���w~v��U�TƦ�O���\�1~�n�WO܇�|�� �]���b�a�����wz|+�)��SU�5d͌���rBv�j slq��W6>�{u���W]:7-�z�˧��`Y���?+ׯ�s������% ˂8؜h����}U�4F�+PY`	�!�8@���Z�Av��2m��v�m�(`e1f�+�qó��e!�>���E��g2��L�"�o����C 8p���������zBB7P���F^A�j�@\��T��W��㾾���VM9:�0}�۵+��6X �`n��=�hf}|�����A9�� �	�u�Q3I�,�L���2?}M��;'ؖf��1N{"�zn?N?fn�_1��ͤsk��[��e�yh�a�!掖6+im�n�e%�r��h�*E�*���S���������<S��W-�$�:�|�����iK���m�<i��O]��c����h���o��an��(��9I�*k�-xk$�Oݯ�"k߉�{f^6�G��Q<Is�t_��daa)�_�&n���)��%��Ce�f�
1+�LBX|�j7X����5���x/���ro�AI>N0�_#t$�^��e�d��h�9K�4�jwd�˵�־O�Y�^�G�����ݏ��g@�jȖ�E\MJZ�D�1��#Ӕ5_0���0�r�+)�3W_��#�ė���Ma�պ��Խ Zp����ʯq�3s�;h8N��ڧ_���^jM�K_�K�>�g�����^C���X��nGOs�G��ߴ�##�%�[H,�5 ��#*X��jn�-L+�-b	��5 ĭU�[�e�N�t~�pu����a3��������S��9Ԥ��f^M����,���s�{�������=�Pꆝ��!��G>�ˆ��'ˀ�3�Ǒ����֐�7f�Pg3ZGU�ȼ�;�I��rS�Mi�v���6NZ���D��St�0_hu���ѳ�E�$UU`��Il�+,Ta�i�Oݯ��jrV��΅?� f�A����h���Ds�:�]���?^U�m_%�6��'��j���D�J��2�(S�%m^P��ommM�l�w�A<x�e�!Lw!�	AP��ypo�b���������%���Z�P��Q|�.��������ހ���P���X������B���0W��o1��vw��",^b7���������K��`�'������K:H,*v������|�Lj�

�b��A�kB�-N�����z]��{���l���\�r�Wuu71I��!L��^�����|��5���d�ǁ�_�������t3���p3@����S�m#ԇ�Č�%fem-~���ԕ���		,T�:��I-)9�-,�/4P� jN޽{����b��A�[�uC��\K[��:�^6_�=2]��������t}c�L<z~�����J79U���10p�^��HO+'���4+%J(�Z��n��h� �'����98$������fj�#I�?}�_����$���������d"�J����r�*()U�����F���w�6dpZ��1g(#�����"1�YIQ�.�f<ʊ���x����-�Z��c���So.31��cG"XF�����,��23���9PʃQGJ�[���uQ�+LBxE���h5���2�no7�s�U���"�yi@�z$2�$�4p����@�O��kt�9&�:\b��4������% �SL��KK�@�`�"��aDEe@dHZ���^q�6�'�>�A���cԶ�|ᒤ�{G� �9��0XlK�^1��y���S��|w}�,`� ��Ԓ�h9�)4t�4UWWo�H��Ͽ"1����{vϊ�8m�i*�L��:�G���%�/f�tl�sO=�Uv�[laBX�V�y�=���gq���|�gĻ�����Ϗ�צ`�M@��u3[�8�u�ˆ/��Uk��hK�{��+��i:+u>�;���YP��!�G��8��D:���<u�ӑ�!bg���AKc�I�H8�#�d1��n������L��V����n�3k�f8R��!�-v���[���`v_�J�*+#Ø��]��bXQ�&~�,�;r�y
�vxm<&b�Oo0�Ix�</�O�@��t�
~����Bf���WP��y�vZЋ�q�-m^k�󻢙�[��
,ڀ�K�~�v�Qh��ȑ8�o��eEa�'�QWW���30���̃N�)�#�MM���d%�x׏q-H�P�����ƍ��_B�kNNW-�����{�S�����AHB��ՔR*uۣ�!
e��$ٝ�u�ܥ�TF[±3�H�Q2Nq
ٙ���}��޿���}|���\��~�����+�~x{K9Y)|k�KQ?5k�܅��y�isV�?DC謷����]p5#���ߢ��[r�&����ƌXo��+��6��G{��5ާ�U]�U�$�O(|��TNR��W}�|�
*eV�Eu�qк��J�
6������c�>�Q)�&�Z��,c��η�E��{!�u����7��ָ���s|�A{{���Wk�X�^44��)4�9ʮ�=L��4�`:�ߊ��ee�#�J�
̹�STӮe��ٴ�uA9#��6'���m�.A��/�߽{W"iq�-�N^�c���e�(t��cǎ�ӥ ';8{Μ�?mqm'j\��`��2K�6��QA@c���n}}�Q�C^DC�
9ή��$���X����c��bh�?�4k�_���k^�~Ԫ��j�ܹ��x�b�)�R+�^�}�f���kĕk�0�b��T}�G��ݷf��@ݪ=|�0VǢ���7-�m���}
p��}@���	�r�#���JVw��d���38lк���IJ�Tg}�=bBY���D�"���R�����[N��0�^��K����_�ɖ�b��~f6.����*�gQx8�VFo(Jua��u̱+ݺd�]`x��Fk���X-���v���<�.&w�`�G��o�x�0�l�*������C������.����߷�*�u�2�B �@pʑ��YbƂG��>��ݝ͖#�܅�5]@ԊP�t�e}hϤ�é%<l�lצ'�T����S.���Vd2�s/�`m��2��v>��	���Y~��P_�sC'�,�>Ύ�]yy0��>�ps�I��r5ڴ�س
�z�"�����[D���?o�&m�d��E�M�.$��W������P�)��C�!_�ti�|���ǻٸ�������|:�m�e%��6����)b���u�h¢�N(�ӎ!y�uKZK0��o���2�^䜀A���ką��KR�7��g��P��W�XNk����7����_�$޸��Q���P7?G�O��S�U�"�|�bo���s�.�1� ������g��l7�$�X��v �u_��1�cϰ��"f�:�\3i���@
u�Fa{7��#x27�{�o:��S{Y%M��)-���h�E���a7_k��Wj��#"f��1�P�0�ƫehn���A,�,*fIQ�]pO�:��^��Õ
�������\�m�ҩ��.&��)�f *����6���{L������j�(��)�1x�ÞW M�]��Z�14���$��L�]�Տ=�	���Wg���)�\���$[���5!>����}��T�{���H�G�o�w8n��V ���3�]#:���L�
ʲ/�)��sG,l���v�-�w���E(�>��
�:1+��i1i�ڽ��)�0#��e*ea%j���F�PI���<��I��A�py���x0�� I� ��v0n(/�0B~�0���w��]��T��q��$>[�,}˯_�^�~����`t�or�'1lo@e]���o��֚{�EA�jG<��G�кyD�xC�Э���1�W�U6|���{8@DxH��z��^�Z��)��D�#e��8"��g���ǂ�O �v�A�Jp�p���C��߲~"B1-s�&$�s����1Nԛ�jԱc�9{	A�M�	�kOySX#��p@��1�������Z�-a�S>��Ç����fϛ?����@��%JC��~�=���{�Σٝ��S�~���A�yL�Rb��̚P)�$%6�ooK)))�XM���߷"�UVN�{��ڋ�X���!q����sj��v^{C��2y���ν]M������/P`l+�������g5_	A6�	B$��u3+p ����͛7I�7�;{�WjFcjw2���O��Q㥵��|�
��0�p�h�}Es/
�P��4���֞`}���ym��	t!��野:9)�g��d���-�|_)GЉ������9�Zѝ	���^����V]=��P�#�~��{k`�&�E�����w��k�[�������i
j��y9�!I �85��R\#��{C�#��<����/��_aq�w`��Ova������]�V���B���:��%���w1 ���lƕKh�(�w��>|���c�֠*G��r�]O TG��$n��PJ�����1��D�wRe�@W'���]���NҚ�s�ss|����5�D8�|���(E �n��������푹m��[\F��:��'�������t|؂��}��r�> �#6� ����A��<�#�f*�!TZ3�O�˛�[֎y��!h���3&&��70p�&��z%%��|��3��b�����H?qiPC"�@���x���R~)8
c��O�Z��wN�����
�O!�����
���������l_>{xG��'�o�H���~�����˟8!�K�[�ϱw=�_�m��Ѭ�U������O�Ƀ2��[�����whi�i�$�D����܀b��H�H�x��Λ��-�%����$���i�M娐s�Kl�ׯ_���y�Pp	0������T��Jt�B"�0�%'��b*�X\�����`���u9��^<D�U���i]|��W���>�=+�~��{�ַ>�PK8T�R8v��@h��́���HSX��zz?�ګ��(U9���p�-Yꎛ��M[Y��PA��V߲�e���jb�p%�4�������=�G)�d8T&QU�!3K�k�oY���v\S[��\A�?몣��]\�o�z�~��������{H	ޏ�{H==k�	>�/��Zk��'��ewg���wk����O�㹗Ɂ�`LQڰ���(E��]��q5x�J���aZ�v�j�*N���(�r�oΜ9�ُ���䙰�Գ���������� `�f����\U�qX%���a��hM�k��<ӒrsͰG^��S�xp�v��֢�LI�8���r�����X�ddd�M�{�"� Q��D	s����w��u�׺)��Z��dI����ᑑJJv ��^�����n��|<;M�N�~kk�C�h�4�����T�1�K�"ܸ�,9}��n)�����L�|c���y|���!�#y޸GӃEe��-.����eQS���*�>���_�4S����i7cc� z�W�B�B�a�V�srZ��@Gg���Ǉ��ƿ� []]�C�k��μ���f�DR���]H����K眓�c��|J��QK/:�d��!+�Z�7��#��.�a�x$�B�LO_���������gdI�Qz�H����N �3/� �d���������d;�sgs�P��S��#�Wd�|� ӳ�ɣ��zt�1)�
� ����>�c���y5��k�����~/B٥��W������y��h�J�W/�(�|'\��Z:�O�!��;��T���a�$�ӍN�۽{7�"ƫ��^WƑ���ـ��:L�����Ş�,f�v�,���w!��Ň��a��a�!1�J8��+W���	�����%�n���ƜG.3��	0Aı�݈����lQ�Q�H�:�hN8�UA��8�����8�c�2Ԛ���!)99����F�X��[�����VI�V��}� �R�o�/0u��Ͽ	^w�"6�)���%�������s�U1�eG@�׸_Xh�����;��?� `f���>�!2<t���{���%��bqɶĚ��(qV�Օ&*�sÎ>�M&`��2����|,�UR�18�,c�
Q�'��czE�Si��F����T��m��+��NK[��P?^9��ԿA#��O�ɸ�v��ɱ�0������w
|"�y�ݿ}[gd�Wd�
��ԓ-s?��2�����c��Q�Ԟ��Ꚛ�ec�8����D�O:��4|O7̣�i���lݍ7����g�
U^��<&�(D�Ȍ�3xE�|�J轧���u���w�n�Y�N�;�N���b��v		%�y��>	�����ێ1��GoH�P�n0'��\w_ {�5c��Kc������:q�<���+�g`�\�;����.�����e�*<���yP�O#�]3� R�D�Y��&ʫ�w�<z��h�����&j1���ߣP�Q������絍9�<�\w7-m/����'&�5P����n�����]��}�ؿ҄I�T[�S�d> ]I^|ꌁ��ͯx�����ח�=������kj:���"��X����� ���[��8��벜����UP}�A�/uu�d����B��Y��gR��|�v��رc���l�������f��N7����w��eZ?=C�{\\��K�Uk�V�O�ݠ�_T���z�;շ[��
x$���	B,��E3��<�h�G���Iz4�w���/*�UP��x����G�_^R+�TRR2_F&�B'T-`T%ޮ$���SY0� �j�9�Zo���V�_��1��_�8S��T$������q7���L�!��Z��x��d�k��b��o��jT���_���E��7�Hϲe˒�O��� +g��[_W���B�U�\��#͔@�.l֞J�n�$�pnV9�K"Nb�g$1�wpk7���+�o��n��|;U�� -7r�m�^8����ܐ�U�_�<��Ao�pރi�I;�l���}�ev�Y�
=��@3���wg|J�[�0i�'��< 㲳����N����S� 2 !��w1�^܂Y9�A�Zw 0�}E�S�&8E���&�B�	1������?n��\�"�y����[��Hv
u[t�v����Ra��@̒�����������������ne�od������ �#Ft��hȃ<�i�X`_>��� u�Mӥ��UU��a ��y���������n?~����a ���,�	�,e�Ii��l6L�Md7��3+t�9`��oϧ^
E5�ST4��N��ō#�oINN�����ms��P����,"��9�����~U	E#K��`dy�%-��ߟc�t�^mQ�Z7o�����L�5�?_s]������ n�H�����J�q�V����O�jtFh3nv�x�e`e��V�����fY{hA��]i�Y��?���N�r}\�������b�K�������%��_�L�o�DZ(˿�X��Fl���3wI 1�'Z�mlR��R��ۯ�$P/�Sx���{ο�/Y���w�|b_k���"�`��*7 �:E��2�{�VF��P��h;���
FH�k��.��I�7:��jɢZC,�ljpF_��,��l0����D�35S!�\�N*�5��9|k"���t� ƭ��j\$s\�9��5�x�����:�?�jHg��&�(�;:&k]K#w�k�`�.đ!�
yn*I�#���n�OI	+;p�R7�7�A�=��w$��Yn޼���שٮM���
�����5p@�х�#�q������ԁ�z�e^6�鱿xF���]��S���Ń��p�3�ED��D�x�pbъ�в}�����{��4��{�,F�|i�֒}�1�<܃K�Z͖����r���A�2��^����׫bO�u
'q ��H�V[�I�����LLHZ$�C4�텃��M&��"&��7��I/�	� �T��:����=�q�����۱s��<9��Y�ƀ���*��3�nPV�ܶ�1H����c�#��a����uV�78��x�Q�6�0;ϒA�����}*c�xy�8h��鿝�ې�v8P��߾�gX��GJ�S'�Kg�g]���U&��N� �ƔÄ��TD#77Wq�s/���nږTa%mU���R,(�" /8�7///I���^n�����o"�
c7�=ź�C{q�#��b�i)�@�>���7��9����wꍰ��ѓ'��x����n��^���d�l��$v\9��څG��Ⱍ��s�dJvӦ�ɥ��u3��JHHX�+�/u���Q�B:��Sq�R��<���Y.e[L�v-q�*��h��v�}J�l��(N� dO��̏���l8�:#�d��m&���)G''#l�㧆��s@��L��/���[����W��BoG1��ټ�Y~����e��m�� ����#I]Lϫ�qߊ�8p�S�L`Rsi�k�������&Q�/��I������%R�؃[���oU�K�oX�z��%w��=R�~��qZ�{43C�+�~ �߿BR$�E���5n�����9\f����V���
�`���\p},���R���ے@�nͷ�@��]���{����4����TW'��vvއQ�Ww?�z:��6h"_��~���n?�ر[�r�~P�J��q� ���,�ދ�0�/�a�E{�s%)��i) <&���bt�y��_T�E�N�?�˾C���>a]��6mZ��J-��?w.;|�i�H�rQ����s�fȦ;�Л�!�� �?g9��sR�����Y��l��"G0�N..�I�]'�[X�wb�8�������k��)\�sj�#�������K��_"�:]D���{�S�j�4p4�D�x6'��~F��߽��W}n�oȣ'O�s���&���:e_�k�0��P�ZW6��$���R'jU��Y�F��Re}��A*]�iˎ]�*�~�ڋ׫�&O����oư��70u�A�>�#�Y�.���VK8�|LD���##�o�5�!���rTT<���\��C�w��[��V����O��Y�*�ѣO��"V��q5��ҳ��#�,�08�r{î��PDS���C��6 �]&+�n_�bE��w`(��i��͛�Q���	�A<mِo�sf�?����)���Wq�(J���y�X|S8���R*5m��r8��<&�~SbLq�Z����;g��mp�?J�����уK���*hL�м�<�1����2p����P��k�iӮn_B����q�+6��Up�E��B�ԯ���^���A�;^��2L���;8쪑7��h��G�֚�t�A�-j;c��֌_�B����F2"S� �imm��R�y�He������W��MI|U"""�{�xܬ�VN�E�W3�u�֍���e7��UUUU�Zv
�KvS��������qtt|O\�`g̷�B�?	����5:]D���c"	_�R�./��)�M�������V���4S�7Uiv��.��#��'��h
7�p.���$�5���X4�6�̖u���%[�,�7�/�9�����Q �V�7��R�S&�S�榟Sk᠐D!!3�L���K2��ʢ��?53 p��B�Wk����}��+���!���X�:=�JM@ta�~b~�N�#�8^�������	�"����u��*+M�1��\ʗǏYN�}��#�h�]1��-�d�_p8|x�\wH�w���jpW�t��̽��n��4M�}J���c���Hn�I2b�p*	(\
���K�(���Z��!�C��10,5jv?~���ym�TI�9��/�ck�*�zX~��#IK[�%��~����Z��N-����T�������??�#)��7E�m�ْ8:��m��*�qFFI�UĨ�TZlS�@xp�$���>�:���o�ĵ.t�S�7��J�V���ݳgO��Lmƚ��.(�h��Ɍmohh�y�fzE���v�C�bQ�*')ۍ����+��u�z@��def���������?z����]q��%+,]�a�^н��-i��Š��ޥ~>L�xePn���o���Z&E�8�8��H8�<}��P�1�ʦ9�$��f=~qS�:���gSF���E*尪��+ĝ����TMC3����x5*mml\*�a�ߦ�$3��E����I��G%b�����\��իW���̳׀jTU���WLu�[P���;��+P��q�>�D��=vLo��f��x<16L���dc��Ң�,����z+N�@h�5�ܙ��!$�6�ب\�����"k<��5�Xg������f��>|�ELߦ�F��βBLn���Ȫ�6^�яHj44>��N�?Mu�$��9�h�ؿ �
�9p����g7a��,������oV��<&o����?l�d��(<"Ű�y�����A�w.��Q������A\��;�d��k�Kaar�!l9&��
d&*�=$uyGGǐ�4e�q2��Z��ÑNg31���v!5�A�^]鹧�*�
����
+��]QQ1.36�e�nG{�WQ��7G��MqXyu��!!Dￃ�ǡ���v�0-�����AL=����9cl0��y��"���T[ԧ��"q��3@i�l�_����R�&�9����5X��%e:E�7!$�%����R?d�s3U��}�@���ȑ�sL�d�-k���
�)##�H�'I���XK�`p��-#0:�J��@���B`%��S.�s�ASp	'!��.g2S��L5$F��s������rq�A+h#E<Μݾ~��ڳ��9���3v�uo����i��.c#E�X1�@��T�g'�D�7YO�R�P�Df�G^^��d1����`��o�
�x�F;�._�|Ϣ��r���	���H������L=E3���p��"Rj�b"�a��ӧ�jCS���K�X()+��x+m8����E$Whq<ۥK��-������9�l_��-�˯b���)`o.;[��&��[���l��Sl'@��'~��3#4�k��&J��uvN�q��.$Ag ��HO9`�@n�޲H��˾��R��N��^%}�,iҩX #S�9����w��Ǌ�+={�^��Ours�:ϳ-�>����3m����k&�����gp��^wCO?�(c� Y�
�	s�$asw�����?���C�UNi�?�<���l�]�neܟ�U{n`����b�O4I�.���>��K�{�n=�81lb7� �h`)�/�_�x�ȑ#�kSl��V��4_D]��:\�G�#ud�W�VEvg�fg�L��,��0>~�>���\\�bh �愵9̑)k����q�j��οd-!�S��94~2����k�*\o�sjCB�3�8yy��L��� + �9�7����,}������Җ̜��*�h�_u��yn���*���6õ������^R&R�~�+`0�O�Lk��t-@�ԥ~���CVM�!(��)�P<䗧U���x���g����&́���Nd G���p�U��ҥKqpf@�sB^�'-��������Q�Zg���^�lq3&�*uj|��X����lSD|4�ߥ�+�O�S���$o����Ȣ.otQ�o��"�JS���[Ha��#j1���"���w������T�}I�,x�Ww�s���H_��A�P ��3�/�i�l�rwɭ��7�oPRR�2����^�c__&^7 $���*޾y�Ъ8�Q��ֆ�?�R���*�vFF$r�*߮��		��/4��dmH�L�#��m�o�ô� :Zw���}�KJI	�<��C��g�p��u;)�V� �]�~
n"p�-��z��_,^|c� �dw����l�h_i����F��f��W�(ܯr$�) R��7qR����p��\<�,^��0��G�*��svN[n/��>env	 ��l^�a :���0G��s��דd.6+`�$7�����|�X��]��=���M���~��YȮ�~��$��5n�n6�":k����D�����WWv�~`V���&�6����t����}8�)Wi��4�`\��,Z7��鈨$��E^�z��S
ov�ThqD������n��Z���*�BG.n��r[��v*u���=��Hm7�����	F�!.��V��t�w�������'��\홨�����]��$u1`>$3�bwm���T�R����z��8�P���RD��zff7HsXĆ[�8�erk����3�V��*�U ��Ѭb9���5JS�`1�V��ņ/��g��U�8�QM��? <'����)ld��*�.�v%xz.�~�h�9o�����M���$�21I����<�c�MNN�*K�� V*ϣ����y��(�e(QD�8��f�Y��2�����W����l]o M#�w?ɟ�Y���҄��u&v� �C�����mb�4H�LR� �[
?*��ҠF*��|���!�	��n$'$�qc�5G0Ŏ �,�颳� ��P�
2y�~��ݗ&GNfzMz���6^>�p׮]��1QQ�]_axr�[Il��s�=�k�&���1 _��#_�g�[YŐ~�𥸃c�~����;d4��S
�"+#��V��7��5If$��,��ǫ�+k�	�-ux��~���{\����X��KC�k�	��g_SOt5�B�>e�֭G��68�J���<�:�hRL��T0�D���k��U�
P�8�ϩ���ځ��3Q&��h��%s(��L�:7�3E񉉻&�	�[33[�l��S�& U"#E
lwx�/��, �r^�b��7�{YZ
2��ؕ	��s�*"���x�=���60 t2��I��o������r��qq�.kh���ܧ��ÙQq=�T����C�i�/�yx^�G��I����w*h$^�o������u���@���p�%�B�'�Ys'����N�D
�F���6�^��7"�Kܟl��g/Δ�}	X�b��Օ���}�aB�����A�����%19�=e|��ӠV��'�	P�^�dՑ�M�M�zx�OVB��Qbbչ�����kr��=�Z���B��q�2����VT����,�Ҧ����܆���̢dF{�'2�zws��%�v��_k*l,�G�[)I��(�=�xV�_��R��&Z�Q�[��<z"��*�1 �0I�Z2��O�zQJG���$p$;0�n���탟�L���o�+%��E��N=h�h�Y�T�W^h+�`߸q��$��f|�vP��[ d`dBg��0��p�T�+bԇ9E�N(L�GbKQuKW��d�*���Gw�0h�|�������0M�14 AQ9��Rd���`7ܸ C��8�	d��
b?Β�jTС�����P3/La��c[E����}�T�䫱�ss&DS6�����(�y�s��`��R���sY)6��1��>K%Jv�x�@��
3�pb�mee���u�By�ͪ]=V�KO��{��32�l,�D�ɒe��Zb���:rǦL'�a��%M�l��֝=p�����3|���a�evM�CǓ��A��C���h9T���H��i��Ƒ����y���t�*Ku�k^@�5�>^Ҙ������G�`a�𠟟%�{�@;�?R�݌�[,kb�y�-F`VI�/��K�ڏw6')�]U����1��J��n*S��=9���~��`uE=��b�>0�G.� k�Q9R��`�\�ȗ1��`����>\q�X�1X{:?s�;�<���bDn_r��QG�r�'J�M%���/��[_�~�W��o��%�גV��)*^�]o��1�.�,��_�H��&���f��%��L��ES���c�iBա 87�������EEI�>�X}}냵dkO4��⼻fF�3��t��?v;�GwLB��F'>h���A��������E$:)��{�HЌ*�E�6+N�(�D}�����pd�����H�tk��ف!����7�@?`���w�y�koGb
	����tRB����)2�1��\��<0N\r�b�>�����M�)&�Tsijjr�#�G��wFtA��-{��`�����.��:C�;)��[w����Ao��p6�5|�>M>��b�ʕy����]�̜A=JNއF������t>�Q�$)Y���E�6���rhI1��z�'6?;���|&���l!��	�/�)�X��Un/��pG��`-g0�8;Oo��/PviY��J2A���EL��*!\o���(c�,�7�/H�� �&+�s6���z��q�%eS��,�H(�ҩ?��v5�LV����hb���S�zh|b�[�X6����ձmkq�I���/�]�ޒf���V�(F6X]2l�|�+p��%s����O�z4ؾ5B�=9I��؁��<��є{�a��CSN�]NHHظ������ �aކ�;��O�����O�G	� b�[�-�7�j�G�s��ҿ/v���U�C/K���ּ\��,�Xu\c�%�t�2�ʘ���5v�I�3@ষ���d�������w	H���`D���sc�g���f"��2�s4�)�-�Q��k��f��c��U~ͼ��sf���V���yx�� k+���鞔�c�������������ӿ<���+��_پ��V���%������Z��>��[ 4��떖��Mȴz�7{#G�2��;w�A�S��9�4��q�8��͍��500`w�������g�כ��O�j��'ߗ��N���}^�������q��u��0p�������>&����M�slw��}���'̦E��.M1�,X`� �C���T���6�@{<����	^�d��vC-���9�g?��6a.��/@�O�?T˻�?�:sۤ[�\�n^�v���lN��śkfm]��Ҕ���Y�M�o���}J�����e����j|����`L�k,U�, ����>>�X*d��M��l�&V���$��vo1u�Մ�SJ�ҥKfr�[$K��u�6��>�|�Ot�s/Yˡm��
��Qpܠ�z�i�_�R��%4�A����i�9O���\3R���^�o�p1���b����^��;�9�p4�G#,��s�H��H�ˣ� }g�d�<�(��ԩk��������vGa������=���J轿�{qbb"I���9�,Yw��ג�i��Q� ��6�4��'P.�	�[$�6i� 
S�1�r��l������I����j�s�T��.�*�g�ϕ��e���&$4�K��)3\�K81T5�'��Q�7����:`g�sD)�ɞ=\[A�,ǂ���6-�n-_��;|�U�XA�0��}���[*�G����CSg�9�Ƕ���b���7�uf��k
An����=~�����(�#8�nx|�썀�<b2���ėؓ�X��(A�/�<FE19�Np$��U��
�T^�C��J�l˽��ѕQw��ws�j����]����([ ��jM��D£�^�G����X��y��HZ�pƃ ��z�3�D��4%���_��$��m�#F��dO�}����2������իX�I��%����T������L���ۻU�y�\}���g���kV��r���#�YG�� NvL���Lq���)�K�����J��?r�ݖ���SI�N����!=l����<ֿ9̑����`�UY�O������-^'�J(����Gˍ�@:�?��	WSQ �-��2��,�.k�l�Xk櫷�?�;uC%���ǭ	7B��s��q��i�6 �0�F	dw���u�X@����,ƙ�\o'��ߏ��/�b	��q{c^e��i*7����t0�GŶ5�&�������盢��y�G�;͏"��5�F�����m���xh'�o��5�ڵk���ac&n;��N6�F����Dع,��E��<�Bo��^�,�����^YY��A#�:��a��}h�l��4���rZ�r��.�P)�؊c^rs?�r�Od�ó�ǿ��N���Q�*�6��#������R��#��4C�N��6w�|������}�s�'/��1�x��j,�F���<��y�l�&}�\���Q�dv��k�� �a���h�.���'�&���t���'�Nq��~��V�p -�_;�0�CKso�FZ���>�-��X~C�(f�y��ݠ�)��B<�(�������Ç��-#�&"��_�+A���ؤL_��P���!	\5����ֆ��_榦������������"�*�QD�f���J���2|��M�Q�|��Ŗ�� 'a�M�~������L4�jđ���C%\�-XKǸ�Mӝ�w7��S�	,��hcP��ǅMw�� ��R���-�-W��0�`g�;y�dI`�X��<{��M����/^�ѥW�<rJy������$����%�דe�-��e�����K�������W�C�.��u��p�ȥ)� 6�N��t��L��?����%��z1*�"�/@��M��b�P�e�ܲ���8K���NU��vxܾ���=�"��GE�S�pN^]�S�#{������Jy	h$4������#��U�������oY&'wU?>YIl&8��Ӥ.�\Rn��[�k�tl����W���j�I����C�ܼ��3j5�;�g�*�7l��Ө� �@�[��X�� 4k�����y������f�`�Wa�f��ɜ�k�R����;7u_�q�}G�c�h����976��J�55}+��8y�n'Ŷ�D��Ri�7\��=�T�)���U�'#�����|�]��-���wP�,3�RV ^�5��4¹z��}}}C�e(�Nl�.,lD�N�����}����m�^y�D�r(eϟ�!��Ͼ�c�p���EzC��|��W0�"~x%�WW���aF���ҿղ7�::�j��'M��ݻ�*���Fkn.|����[lfh�h}��1�X��kr�&|]�����!b$�vEqZǪ�Y3r5�Q�Ȗf��| ��h"@� '� �a2W�4�W�K�jȯ%_$�mQp]�`� �\��b��j��S]Y��m`Qǿd:F��X7��u��,���w��dy�����qW��+mҸ��	H-��f<9o�Ök.�-k:���3��b�h��k�����Y;�*2�N�pi��c����We8l4i\A�I#A�K�b�P`?|��E'�c��o~򽟅K���*]@���U=����E��`Y�4�Qb��J�ڸ�**\?���?Hz����c�Y��*!
+M�t���沈�>�=6֢�^�6��&b���'���Y�?��t�58Ї�LO�l�����Ʉ�Q����hH{����!������������)�	�V5�%0ؒ]Q�O�E���Y*�>�Q�e�R���Wj��)�FxaV�콆��}��kg*`���т�XM a�e�KǭS�%K�9EC�E�k��'>�Hn)w`� ��Cf��O���%�����,S8j7yQ �q{�R�a �^�~^p�"��ǭ]��� p�~�����Y���J��#���)�Mi���WK�c����J=C��x����Į��u!���+C��!j]�s��/�c�Aw�J����E7v�={vrU߻I��.Z��ܫ�'9'�S*b��\K��ċrsU�Μ�>s���ԻLm�<a�|JXcp������ _Z�b1H��M����l�d���ܠX�����ݨ�{9y-��L2rV9!!a�$A.[��˼_�^а���5�ϡΔ���M1v�,��'dI�w�Y��gX7֬=~o�_�$T��=�$e�	 ����Ä�y�Y�88���O�:�	��׫�.סc��^.p���wp� 7O)����t�Ti���i�j�6�5�ˋ�X��;�m�y�(�Ȇ���/ �:C�[~E�t��!�r��Mar��.[���}���,�����S�bh�%�u� ax:��L�R�}W���o"��t��6��<o��jԭv?�'�Q�f��@ ���<�Y�0��k�!y�B�uS���Ar�k�����&�>�p�h��{�8�鹽�|�E�|g�J�z��c�g����~�;�i�p����3w}�-0^�#w�ԐG�ݿ~��6,W��~ɲ�c�x{�c2��u��I<	e�'�  ��%a~&ۺ'�i<	x���{Zv$3���۱����c���`jii�� �Lw�zaQQ��1��yY"e����Fnr�,W �T12�~�<$$�����Wqq�+ۗd���~�`)h���rI^�����e�	�Fv��8�c���8חp��d�!��1Yx[Cќ<8�ŀ��l.�z����5kn��ԡ�Œ��7o.�]o�B��h;�2E��,ȉ�j��}^b�*'����7�2<O���:{vʪի����h�Û)�2I�`��Z�Zno�zo���E��^w$ڌ��b��\���ڬ�,d5����n��Ӻ[_����Jh��n�ٵ�,ܜx���)��Fl����V9���ٽ�;`h
������Y둒�����C^T����_��v�J����<\��up2��XU_Of	�M e}��̰z8����d���T�H��/.�����Z���Y�z�|��X�72��zt���4���8)	���?޾���rJ�b�`��G.�Yy��wv���/�t���鹩�Q�8�̱��n�Dr������1$�b\?�n���8	
�]�[��Ʀr��M�l��/Ԛ�y��}7����s�T��F����~`B����d-�fג���@�W�J�ұ�"�����f�n�Lڋd����{�HYn�����ϱ��S�z��U����ĺ`*����M$� H+u�1?���J���X��<��)�|S���
'���--���뷹g������m��v�c�!S�$�z�9�RP@K�|��Յ�<�j�1�M�)Sf,AgFrhG��+�'4�Ө�` ��\�톍�?f�=/q�_�v\9X4@����gb�'~��1c'�D�y{K9�ɓ� �X ��ё=O(R�����������<}��f�x���OFQ�P9;�	���|�4� ���_��@ON��|*v�e��n`na1�R�G����ݢݳ�޸�Q$���˿�s��`��Vx%�!8��F��ӑ#d��>/ž�v2�('��Q�&{4�p&��:�����,�\�&b՗� �*�M�R�Yb" �U>�������r�)�E� ���5���ԦdW��0!�C0�����O��>+n��M���p��!v�N\0l١��n���okV��U4[�˒O�[�e��w� #� ���d7_.�����_�E����HxP�]��5x���qs��ûb$x�G�a; e��	 Y?����F]�G�eQ�5��f�pT>V9�yZ����y�����<��
��D�0�UB%U�"���u��y�n��i� ����Θ��[��t���Ì#���3����#؈����i2����~�tb�L�9)�m���*���L���Glo�L�kx���֨��&$��t�0E����KR=���5{�(M�>��EE���Xc�g�;���Ȁ]���O�m/XV>=Q�����6��B��fKHx~�G1r;:�fe��N����P�N��W0�N/�;���������I��d��T�� �͓��z��HQK*{3sr0Uɺ	�y���t� ���6�t��z�og�n�q�Ek��	�Vu �Pp���t|�b]�0I��
�oG���45�����e�����P5A��E���]�5��%�[":^ی�s�䷹A��	��U������jf��������K�V gĵ��p����I��w+W�4��S��~�e�¹m �
�I=�m��f�U������5����38�>�`oO�ɳ��_:X��R�>�t^J�,`0��I���>��M��4���S2e��#�*ob|d���R*( ��X�����?^vl����d�|�Α�����a5G��0:�����{�����8�jժI��v��jf���Y��w��o-�&��>+�����Sj��a))��		k�@W
p�F�������/�)'��{����0v��V��N�zu�{o��F%�@B��&F/��C�a�����c�R�^�p����m��ͺ��途�M���ej��x[ �b8��Г
�p�?�����Hn�@����ؒ�:r���������Q�9C�e�ԯ�T	�����@g��qZ�bk[�����/�����c������䴴��	�i3����6��}�J��x�(``�YV��V�z���K�<<>�Ѿ�X�v+7d�5L��� �x~˦�*�R�7�T�p���� ҵ�
�(�{���P���W-@8U����;�_رt���:��^�b&~wv�I�pϯ
�di�</y��ԋ:����Xٻ���:Ś8���<�M) �BK��)Ƅ;Ǖ�%^��}���fj�@��jW/_�n�ח��-반�dbuT$3Er��r�C=Yy4V��+z��^t���TlR��V���[tq��	����{]������D�p��>=�S���"�i�l��u����K2��۠F�I��O�B�������O�$��ێ\�r��`16ܺ~]Z�'������j�3�����-�٭�ypj�8�N�+?E2��x��K��ȼ~~���'V	N-f�Q��:�C���;)1��Q��(B}�vX ��6w�;-Y�6�П$�h茂Fk�{�*g��Z��Y�w������/E��hL�6�m�y���	l��M�P���4}�E\�=�>yhVV15�Q��M���_�T�V����$�X�|���Gܖ��2�b'�}ۏ�k�0��k � ֈ��g^	y��N��G'����糆[��H�%�)�kee��k�wMQ��)%��7�ܣu\�������(�|p;��q�(�&��I�NpU�Y�|�ʛqd����O�Z�5\���R^~���gEʗO����@����r�ͧ�B��<k�n�����.�LRg�ٵ,���:�*��t
�m�p7����G�U�RX��c��k-:Y�ߒ�D:�Dl��~�Z�)��)����<oџ�giοd�X��I=;`����vh�4���1�0X|��uu��g�9 �-�����VL�s�B��vE~����!;N���m㎿Z�����9�zNN��Z�֑�L��kU�O,`���h/�.;��Y��9�&c=qC^���b��W-��>����Ut�_�3��k��s-��bn�mz	~S�{���:ׁ�:�)LO?h�K���H2U�N�c�2n����[�׉����Y�8W���f����`���Kȓn(��b�u�~��<
ᚸl0q�]5�Z���Ʀߖ�k�����=�}xp���o4��J��;#��{���D?�lϞ�1�^�}7ѺN?N����\��i�k�3`T���4C������<�=���E1�0�O�Q_��}Zp�+p�!��<)��c�M`�F�X�n���Y_�����﮻�;��]�W>�����yt�b�_�<�XSa����H�����$���	��O�Ĩ����Tw�JH���-� �_�
xBo�n39Y�SO�E��v8�k,LMU�R�������U:Kf�%�$�ޜ}|̸�%���x�~�1@$� �L&3����mOhs9��OAR>��������aFV;������Z����'.7���o_
��<DQ��ݨn�jz|��6	�������*~���F7�og�y7�r�'i<��~W���_�^v����l�O��IN<$��B`\��5�C���W�?��!!w���H3ۡ26�jX�R�3`tdc�eR]LYH6�+��f���w<��'��x�������`�S�Ŝ*�M�}e�ø"ϕƛ�ɱ���h?1��w�D���zò����**w���'P���pu۴��c-�G�E��T���2�>V(q-t��ݷ��Eep�.v�Hw��A�<OL9"�o��ג��K����tl������x����B�[��|�ζK\�̳(F�����Y�B���t���U+��ˉ��"����ן�$���p��o����kF���\2Sb�#�E����,��\{�TZ4#�!/�3M����ɒ��]�qL��3A���G�-ɽ�ys����@
�e�w��WǒbmY��^�����G���Y�w��{0�,wG��$��~�(��=3c@���<=�A�=�?��<����!)S��RT�CN�&"s����!�I�+˔9�2��sR$q�yʔy�k�t?�����>��{������k=����k��Y�UC�0C�Y��1�Z�Lz�5����c�eY�k7�g�l�1��͍��h-�)-=}��ī��鰲TTT�t�x��$ëW����7��	��>J�$�����ʹ4��H���B�m	�G�u}=�㋒�9��*�O�Э��� -��~\�����(ڷ�f�A�<���H���H�\ܲ�A;lE�V�w�=Rʍ2t�R�1����iɉ�Fم�/�0�>�&~�!=�9���R? AO�w�fD�Qu�hg����=Z# z�������f�F��<���F��ю�����S!nT�kV���5�'ЭuXp��ڈ��Jن��٨]���Ơ�q�}��Mssag~�@��T*��*����]5����82�5�$j��`��&#ŬzE�8ަ�4��'�ll*�v�ȥ���:>7��+%5U`��wy+*fyp��Yk����^6��CO_)W~׽>�]
�2[�k�a��V�P��雝o?�ϯ�W��V��n�jL���A=�����S����ޖ�Ɍ�)P���٪�l�Bq�OB�7)�.��W���<O!-�"����3�4��MC�p Gf0٤()׫܋�4�l�8�<�hT*���<�XCt���?�{MA%�j���֡�ZS�VYY����}h�vط�h�&)��ԇ;��x~�>H�hb@ͫ�Fn�H�n��(���_3"��dMh�%�9¬	�OGu���0�2�͈}�%`�~��>��=W�3�H}�0���b_��^�r�28�ۧ�ԭ�2,c� ��^T�ç��K���%��+��Dl�.qn(���'&$��3���gn���H<u��f�Ir�1�C=��5773�_FDAp�?@P/Y#�03߁�}ԟnj�|�d������Ν�>%������E<Ǐ��A�f���ͅ�g&�QC�����g���l9<�B��d^�|�ֲkoo����B��8v���w�~g��޿S��}�*O�nYZ>]���e��@� X`5����-c2"8x7D��O0i��Y.Ȥ��zʷ�F���*5Hy�4\4��+�7��Wf%U�h�������g�=^lEm�ۦ�ɾ>���-�tNpm�l����dQi�t�!�eo�E��?�2�*��
��68���V��[ }���D�\�ׂ�v�|��čL�Ծz�e5�YQ�M��(�(�� v�'�
���ItTH��'��~��-r���{��(����>q1A���������0���⒦clE�c�<��;�h0�7o��bW������<��B@��p��H]�F��C��/��R��� �6;��.�]V�Kt���R*���|�.K�E��t���/�e�aFWOFh��Եn9 )̚��p��,+K�u���uvC�ͣ��9n�'E���"���!z%W�-!�*��pk���0����+���5�n�G���7-��ǩ��9��y9�l�ERJ`#�S}�ml��5~��Ѭ#���ASPP��oK��U�5�.϶\+�]"���#jFE٫�~�6ȅ}in���i��WWW�ܥ��Y!�A�j\��t�`�8fDP&>']�Em0�ֿ�O�MI��6�B�%�Ȱ����S�S���� ������������N�z���AZ�t�����s\��67��{d�*>�7pp��$��hI��3!������Ri�nf2 �%���@�6S@�\d��ᄾv8��ތf�H)�߿����HY���(?=Uw��djM`��DDG���3��u�-���~0xIxX�]�"P�>Ѓ^��[66a�I�~�\9*��jZ�ͬ溂Jr�V�	��ب^�w��vs��$�qskRC��S���y������֭�232Ӓ�ǐo����1[�t휉��r6�%�����Hrňmh�S�����}��@����S�Қ��4��=�Cjk�&˩���W��S`��1���lHvF��=���8D����]^vQVQ1�7�I~	6&�����O�	X���y�.�}�U-&�*�K��i�:��&�5��Jĩ���Uj,�.=�{A���L���l�Ȭ����pWF�QQD���ׯ������r2�T�˯��Vwu-�K12�ʳj�J"�!^���S$G�.<�6��(�y�tXx�������V�&b����� �n^�Ì�h�^V�46�Es���G� �̣,5_����=�<�"
����������'U7�v�w�̙�xb�X�U޾|����c���PaxLPP�ݽAib���G:�:\f���@2k��ai�1Îl�>��������?[H��
\���^1�i��>R29��� P��i�^�I�FSb�9)����M�g@�[=�TPm�.�ͦ �_��7i��UcE ~ڟh�R�no�Bs&G����vH������g�IK���]=]�顩��
�H$���ڜmP�TW_��XM�2���z�܈^�ׯ���Nѳ��h%�z��Y^Y(,]V�i���:%ƃ��ƽ�Z��������H��ZZrF�	����W1����D�;M����s�������LL��eb���}��$ ü/
 ���O)[���Ol۳ck�{��˹������RAS����v�\�t���2#t�{q-0C�9��������%ɥM��]μX?�1P6��n�矱�<$�yd�p6�� *��0�"1 ��J�/zܻ���f/pM4�&(O̦3u������������	i��S)����/�ÿ����;�?<��
a�b��I�N�����a��O.�C�=
�y �f��G��"�>Ӽ�t����n�G |���,�.)����Tj�����Z�3�_��p0�uv���=�E��< �:�ux����S����=z������S����-i�=�S���?��Y��LDcEܧ�����M�����e��y[:tVX�P�n�#�}YlF<�����uZ�~m���h�z'E-������oc���H*,,|Z���F��&С�͛�7Yo@g�
{�}���4[~��|Ւ@���ݻSO���8��v���G���������o~H��v�43z"1�
3U"D����\�e�4p�tԾt;;*���ʐf,n�n�\k���~my��sk~*uMomm�;Y! �iز�|�d{.��A�����I����ȝ����`1x�T��v%�<����B�m����^pv%Ӥ���c<x5gimoi׃8^;��HO�v��=��'pp�����r�`��DlI}},�����m�`Uo����Xs�o�w���>̏H6pY���<�¶�����`5ɪ��*��[�'�
	~��o1	hmjJ��X�l2A&�s�����{���GϷ0d��^�Mxn,���
�K�����`�~�v�D�5_�j`ڹ�����j��ܠЌkp#�.'Nܭr�g,BeL���pq`f�S���MWT�B2�p�V�ޏ۷�װ5̌�sHd-5:�&�
o�y>��f��G��8\8*7�z�t7�Uz�?�v��
����ą�jFN�z���GC2T�qh��bT�,(�@��dl/z;3�D����I�����xT���jo����|0k�eB4������n���t��<-��s�o��4��a��Z�XW!�O�����a�Q<����m��)���ͩ{��U+��99Z�+w>qe �C�i��Txtt��ľ�M�+���ɪ�b�T���RBZUUU�=B�;#�y�e�54pD{�ӽ&l���t:'�.7g��@�`����55�d�����4��s�`T�}#�9��%?�5>��?��(V�G�@nYǲ�.Y�(}@'"����.w����*�0*�����5�ǽ��ph��V�d����\�!چ�h^-���7~nGXl�PyIQ�^�J������V��_���gt�w�3�g�Z|<�#�7Ղ�MIN�L�V(�s&��j韃�sO.�H8�O��6Q���/��9`-䢮5kXW�h�3ⷸ��+9s��)��H��S�K�˗����2��������}Β�?���V`��4[l�p��@Z�3W�@(Z�9ֺ�:mwJ���N���ML�8;����HAt�<��4�n�F������b��m�̏KҋJW���n�˺22M�?m��͎爠����dr�A�Ï��[��׷�=w��w/�o?����B�����r�����X\v�f���ʥ��n>/���t���/6Bd�����Ֆ�7�==s����?d���\�I���-��1eU�a_ -�!a��jf�VC�%����G.�](9�yƣ��S�{��0���ں��E��wxy4��W�f��O���#Eed��<�����A�!ת��s�8'D�'OhAzZ���
�ۺu+r���CF-p�������V�YULLo��:6�j��l˞]"��`7<���#���H��]LNL|	�����i;~�x�x�Pn��)Njl���b�Dw;;�xS+��{MF#� �h�al��@{]z��y�Bt֓lh��>���0���y�׊��tP���ވ/�sJ2�I���x�jC35��������^��7tCa딪���$N�v�4b��l��צ�72��1��A�����S���.]cz�]z=�_�LMI��C�愊'��cd"�q�3�'��Z��;�GӋ�GҋƟD|6~����Y�A4���%K��o9�c?��;m��ff��Y�ݬ(���W�B���9������?��!M/�?%vQ8Dq�[��,+=���Η���v� ����ơ�d􀓥e
�����V��*�,M��F*˟�{T�ww�Z�L.�B��o�q.�,��>�Y�[��gf��×��/&����z�x�d_nϔ�y����4ؓ'�δ���q��ZY޼)7���A��dՖtK��
5;]'���	����3,�.$����ʷ��(�tsm�"�c��S�O8]0D{Z�FS��}ux��{[[�7�z�0�'��x�[�x�Jn�VjK���n=�ٱ|r׾G�ׯ����E�����RC>����׀���I�/L�Q�3=����I��\����~�H�A��U��J�|��ti0RSx�x��ϊD�pP��g� ��6�36�N��Yn�Y�Ҥ��Ł��Z_�9�J�?eSP ߝ��<Q�]���Uk��X}L~���	稞���
z���*�����R�=�����c��.�n U��@ܗ�511I2a
)-��D�ſ��*�U!������RZ�_�a����-X����'��:���M��`�)agZii�U��9�����f+�K?�YRt��ԽZ)�]��$+k���H�$z��Pij��aw|g~X0�~�V�p���-����q(\@dN��d;�yW�=���U8�{{S�v��-	ԝ��ɹ��S�šR|��ӧ����=�)�F]����K7H0t�9���}�g����OF���0 M�\�b�F�LtR�1��(�w[��hT�1��zN�M{I��>DDEs�o�8O���/033��8ZBGGGGG���CBn#� <�]n5T1�ɷ
�
��O}'0�r�Bj�6�^�)��֋	�]-����>"�(�rJ��l999�p?�
�5}��1e��f�TGѝ	��*�p�u� �d�S�����?h� N�ם�$834��(�n��l�61�+��x_^�=W��j��f�1�v0<�����r��������ۗ/?�G5vu�(1�z ����$��^�kʵjsNC������~}Ff�ߝ���Q~}�]��X��;lff�����=n���^�u�G�8��"���p���9�V�k���7}G+�3<�$�~�j�H�ش�}2:������&�25��Db����_�����ػ�h�ILL�U���/��(`?���;%&�S',=]�t�_iY�*jC 7'�����<9�?:��a��I��D��vg�P�d'j��${�� ��\Ȉ���#j:�D��(vxXt�f���j��O�6?J:�I��P�\�
$�Y[.G�:?�4�|�;6`/�Ak66d��dy��l���\��t$&��0lZ���g�"l�ݸ9P�8Hհݱ��\,��w��r�;>ӌH��	VVi��q 7S���Fuxn��W\���B��\�P��  ���}���cy�@�(�~3�1mC�j�� G����C���~$T�S���[�i3Z���@ks�H��^����d����HҘ-��qk�>ڥ���&Z�~F὿8�������^�V��z���EtL���D�!*`$I?9-=��{��ʑb��9���N�W����Z���*�MF�����0�Et������Z ?ڋ��Bt+>���3j�7�T�w7
��k+`�z�_*w�v�����N���#@�Q��W?��#�2˻�,�1�CCC��$�Q��,���Q��MWEϰ�/�}�s����90�Su��n�0+uC�@R��O��O�<f���$O�vN��^t��X�-�:Y��=������K0���[��T40�(==�cwS@H���;��RA�KF�����"�{�Tt�����4�M������Ӏ�H5&��?ʆ��Ӓ��;�� |0C��C�}�]�rȆ�Z���!>@���v�1��3N/�)R/��a���7�V&N@���L�F�@���=)d�c��^q�����/Jw��ް�����7^����rrr�З�M�����,>+.���vp\�$_B� �I-�υp^���꤉;m �4�x��dnv�håÒ���=�J`�;�~i�'���vG����UD��|����.%"�	�K}��6x"�n������@� �Ъ����C:'�P�"V,( ���v`26x��w����� ��/5.��nu���3��S�K��{���Wu��NZ�xk� P��{�AV�I��8����<�	���k�5[~���Nq����ɿ|y�}����l���y �i (��V��d���pO"���C:��c5t�緄`���*��C�u�����M�����\����n|N��7Ďi�P~z1���ԢWI���ǃJPVUE�xЛV72��x��Z��ٸC�//������O������}s�@�=p�w�:JJr�j���{�Ym)s]Or_��k�n�=�0�����sY��� _�L�If.L�@�M¹��ׯ�p���D�5�3q񒅒	QNj��ZS���l�)�[�e˂^׆���UIa!e,������0�`�� ���=�.�^��' q��JN�sn����B	��_���p�PÌP��I���rWY�����B�Au�̠��N�B$������:�B�c������-�p���4�b~)�7���gSRR�lF��t�MGaN�F*�"���(�A��˴�L���&��o���A���Cf�";0~���ʷ��"�	qZW���&t�O(��S`�n���r�
��jLR�T����c{���u[n�T��%ي��^gh����yD,q46�EM� ��C9��#
	n�=��E�p��#+�7b�)R�l��������K81,�KCC$8��የ�cy]���3I	�$���4atc��-t�y@�ҝJ���[XZ6���tU�Rp݃�jOV ��;xw뮿�:��ݫ#`N�p,=�F����=Q:�9��C�}RSAa�v133+e�� 8��������3�0(r^��,��RK4 ������ǫ]��Ze�}��'��<s�I��0<1a�]a���'d�5�<�<z�X�%�給L�[���M���Ma^`+��������@�[M�e�!�w>������"���¢��NF�����o%y�.�i��^t�{�b�C `qT�`؝��Sz6.�^X�/�������5 �{��7���ϟ2,--�������VQP�5��dw�Y8\�eG$Ľ���|���d<s��ei�ث4���Qi��p��9yy885n{t��m�G㫹\�P���N�n�D��{�*�S*�[�1��3������AΆҗ�41�����׀��eI݌��FȊ�{�,`?�&
]@����K�(yV���D��;�ӿ>��⢥�y�ظ��WKSS%���v_3�m蹖�����Qg;y��7#'��h�-ϬP�pB����2�g~U�v���b�j,z�.�<�ͤߠ�Ĩ�`j�а���^L!��+�QVz�9����b�Z(W�'"@�d���	�&��04��׃q�ʠ�y��W�y��]pf��i��ojD�:!Z����2���s�\Z���?JM��lkK���.�
8�(���� �C��a��1��t1�>5v��R�����ݫ��|�@�RS���	}�'�(6�߇�}3���N:�����p��V�������JsZ�`cg?�I��Ã�d7�-��Ey��F���W���
hp�01�춃�&z*.�9�h�<��A:�rx,�3���ֿ{qim�+v��V�H>����%e�z�r}Ij,U��V�j~%��L8lj�/P�h��F��2_�j��D;�s�c��̨���/f	aZ�dVt����\ZA��dD�j�7�r(���O>�&����;��|�����T�(ZR r�4��8�j��r��)R��g]pѩ�=o1�FGO��I&�[X(����6���-ԯ����#�?_��&��E�qCC�67E�M��.%��꾺GN�4g�����Jb�b�'kE9�O x�� BO�����ٔ ���&���G���u�n�;��'>/���T�����R(_/4qق��:`H︂.�?�0�d�vZ�D���:�l�a6��MC
���#�c88 �#�}/���x96H-}����Q^�\q3]���ato���$`�"��́\�ޏ>�%�w�<���﹒2��Ǐ��G���qm�Q��ؐ�����Yt���@���o�V�g�Cٱk��M;�Ԇ!�[(K6�⤓eTVQɪ:�I5�lc3�n]�IIi�}Ɨ���"����۷o�yQ/ߑ��0v��7�u��zt��:�~��Y|m�ݰ`��8$��w�ײ�Ǒo��q[|'�}��kq넑z�?��K*ƚ\+t�/Z%�Ky\kk�'�e�!�7�
굼��1�E%w�lM���[2�\�_�ݕ�^o|�)(T�c�Y4J�g/��Ѝ�\��l��*�@@�'� �����O��0Oɕ?�.C�޳S� �x�� E���r� %4�����$����񒒒�aς$���m|��y�4�y��O�}��4�J���m������_ge}���p.���z�D��{�ǒ�4 b�'#~���
Ľ���-[������߾����K����/��N��0�K�v�������=d���rl��<l���en���k��p�����Ν��F��ʣ�����i]��*9��ڵk@n��g>:�_�LDTJ*Џ�B��і;��4���2�b�f�\~�]��뫫D�a-P �8�
J���'ڞdz�O/�p�bMY�4��p��aVz�{�~��V�[��x�å+�&�{iUNs
�o�M�'i.B鸺x�Q�uQ���Io�����U^N'�*{���q��%0����:Uf_��*r�i�����.Ŧ�������m�\őc�L�>��/rṔ��?�2M��E�,(�����S�:ι]6�.��^#��aVR
�"U%eeF@�?��l~1궀V��C��)=:p��$K7�W���|��@������=j$BQe˫�t!B̀K��K�%z�����(`H���b��][Y�Y�!�f[Et�\��L̦�xd\�8��r��DW�)����v�����ѭ0� cP��
7G��
��Pޏn�疝�x�~:�;�ݺu�Ng϶-��0~��)>�F�M�=��3��*Mw�>��2v E�qx+��+JIIYMݱc��Qcr9�ɀӓg�^S;5�8Nne�WR��z��SƆ����'%f���H�e[��2YA���{��������[%F�6��nߪ���2^��oj�w GН#��\���(H�ķB��>Y�D�yk��P33�6��t�f�_�(Lw�� �����N222r�w�,�?+��o��U�qO�����-?Y}�??aH'=��y��X����{؎11�vHαm:Ha��R���DͣU��w��t۲<`1�Yl\��Q��0,tB/V�s���F����cS�W���Y'�����v�]��uN�;��S,���h�:u
�O
��޽p<���Q/4��V�9Ǆ5��=�oDl�bfU��פ�-���
�(gB��Z�k�� ����b��*A�D��>�/�H�q3#'��'�� ��tC�ǭ!Τ�,��[[�������ck�^���n&���	��˾�����4waAa!!V�<tL��X�U���,����F�����(�T*�L����x��Ett��]m�{��7o���r1=-M�A5�r��U�`v����f|�n����,�����纺��GS��F۲s�H^�`BG;nY� ̎��Pcn��gC2�.�w�K�9��D+�z;�ŋ��Ū\+�q~E�hb��6O�V�i�P�1��Y�� y%�̏s�}�)^�`�4O��mq�e�������$�Sy�ad�p��CE?e
̸\f�RO(v�t�h���W� 㱼�&�IQ�04\��nh�u���D���ji?�e� 	Y}'�G߿nq�[���iAAA�Ƨ��p��N�(+���G�ڬ�����p6D-���+X�)`����Mk�?��Ս ӾJLK㜛�#���#�ϗOPݧ���uݫ-��`�|�ܰV��]����>��m�$`�F�%�kc6)���8L�(���U�G�n��c�_r��~�v�9�R�=���Z��KhF��޹#ٗ	��i��ߨ��*d�.y���^�
��U�Ⱥ�;��>�42���c����Y�fQ�0�_���ܻ��a�����7�!�Y��BF��LZA���1L1/�f�n:,*.�1��Z ��Rr4�cx��f�7˰ә��&)X���w̎��5�����ꊉo9*dY0D�a��Q���|�=|Y��Ff�l��;������J4��p?P�JCJq:D''4�(�����^@��9����}r��p\���� Sݖ�;�t<+ �Q��#Q1 �Mŀa�]�T�6߆�]��^Z��� 5�����S���R�t�5뢯��'���Ad+!({�LA��՘�{'#4AFgyN_��\�(�Tb�+gm]���z:<��N��@�<�������ì���K�#�,b�\�dVk^�bB`4���!�I G��h��˖������a1��5&��d:&2�����VDo����8���8�՜��y�T`��V�!fH��M�B�?�;�����P`���<�<�`��/^�@�>g��sph��x���'��'���.s��Ku���n���gv� ���s�L�H�ޚv��g�tu-B����G���n��h��j�?��XJ����<�T�"��L�gb?�݁sE`:w{�W���y��s�DMCCkm������Ӄ' �����Pnt5��X�$#��D�@w����/x�hi��i� R�˝� \�԰�������hJٱ��O
֭��t�J���z� )�ItS\�[ ��B�U��������5K��[�g��mm�g��}2�^��F�� ����B#�M@L�$&�(�k@�(ˣJ���a���N�:s�d|�R���u�M/DOz}��[y���j�L�t�E����e` �AI�[�.��\�=HZ����1�K@mP��Uvn��]��]��m|�fg�x&�N��M����*�]�"��㉊2y�v���9�YMwi���n���9P�����%����N5���zD˛�S8�T8��f2y���	%`����s�����$�*�|o�vY\��)��OZ	â�jj��F���Sd�3Am�P�1���j%�#�o4�+�t�M�[�	:RC%��e[����IK+.a6�&C�k�5a��`�w�Sdy�y���{�`nⵒ�eIY�@&�\�&++���Q�F)B{��YNW���{�jF�ƋI	���� ��5)���w�ڟ�nsS�}��Jw7�	�,gF� �]z����j��K%q�%�[YXX����ȎsH���m��agc������4i5����>�����A������:��gx�o=d����#���au]�}�#�u$���
t�*8�O�w��|�8�v��5�n���W�DI��v� pB�7���z��˯#V����w�v�(��IU� �Q�����b3}Ş��6HЍo:r#,�>L���e�)$��*E�"ܯP6oyֈn|�����-O����q:Q�ş������[H�Ot��/>,e�)v]�k��8q D��01��=^}�7O��x%&┰Cs��i���F��{����P��xj�<�G�b�s�d���-�X͔�������$fp���ā'��a$��_��ӆ�Y�+�Mc�B�/�ւ�9KƬlNqV9����K�m����V�Ϳ�4�[s3��k�۷@��>��� �#u[�V�-,-�!'~�T�A�D&�|��_�>�G$q�GwwN|I���ʑ"*Uc�虾��ُ{Tqn��#�@�7�m��o&���Ͷ*��4���T���zRu㘴g�	 �zb��ӝ���zk�d�"3���	��zTD�[��q� ��G��/�����9Z��B���s9��D6�H����G�U��h5.!���4젧Bo*2"�D��)2�>���6��U���p��?�������͂II�sxZLnoO�K�������zY������/�Q΁����j'#D8�o�@R|ܹ����yGeU�c�j��**΢��c:"C`�\�b�BL��F�P/Xf��
F��/�p�گ��� ua���#�k��� 9���\'\����l�!
��>ut4��	�I���ׯ�^bj#zP�L7��^��	'֗���K�Y�"4���_oz�@t�����N�����3��˽sU����������X�z����_���Ko���3X��d}2���6V�l[�@�=fvDXX��)/)9�>
��UI.me�O(FCs?gx�g��{ɥ���g��{����?�x����!/?�5�u�Y���I�!�1ӡ������]������ZZ��o}Tٓ--s��%�7+od�|bPq��~2���2U�g'�ٲU��<tLz��LI@%5�����QE蝙��qU]=̈́B,$�3����N��b�����@aֱ�.�oU�&{{FR�f�4�F���eBB_���R�g�]P&���{��+�o߾��V�a��DY�tj��fdz���Y����J���z�z~Dٿ)�m6z�M���2�Ӫ�yQZݿ/U��+�ɵ�b+_{��t�)��kR��>���D�zk�R@�����7咵F�Qt��t[(-ll�q���gB�[�ӢgӼ�����B�%��d�M>^Pl�(A'[��X_�"�o�2��}��?*�� �ٙbf���â�!��9����e�_�J&����V$,uQ���\�?~��t��1����pfn�O��ɿ�ݔd����F7���3E���۱��������(��4^qμnB$1����l�X@�Z�!�R� �u���*5a7�	�B�	ضm��8FC*v�R⌑�G��џb`�H��nB�c����
|qa���:����{���0ڂu��{�������m���n��463�G�9����o��F��T�g��ǴJ�P��j�j����5����ڴ��o���	����ۣ9幼>Ž���͟�̿�ݨZN[�}��B�:mYQ���9�`��P�}MP�ߝ��}�n��G�wĈv<}�:G`k>գ���]��ڶ����?H;>�	%����~�͒�p||<����F%��5X:	���Ę�?���h y��[���,=�7������')����Ӫ��0����~
�8�j�#��/�Q](R��w����T��� *�-��w�E#�===KJJ�����ph����Z[%�n��n<�v.X��3)���M�##؇��Y6���D�Xc��c��-�a*�y�z���ܣXM	2��/a�v1��,����o���OPb<�=n�P���"T8���j���LDC�$�Y���,)�<S�^���)]��̻����cn���3�M1��0��>��D���K]*����Pc@ 쥲#��6��KI�T�X�L��C��;�'%mj�cv�e�B����?0O��F�X�t���,O\cc㏕΅ҍv`m;�f��1�eKF���������XB��m��gW1ٳ`�&��o;'���T��=�&{2Br��`�4c���Dg	3��i�I�^^-+N�&�ǧE/)0�fԾx�u;_�z칗�t��jsk�0(�����9��t����d��i^��ji8a�Ҟ)�:�v��o�AG���%F�B�Yt���`��MB��ј�#����� ]z�%�(�V�aEˇ8�`ʯKV���� yw�X~�%M@@�ki=� �z\\�կ�݋ε�����t\���8	�Z�qx���Ǿ�ceLf5�l9�FIYyL�+��N��Q�D�1	fv�ر+ 6�+��#�AH�YK*7���띉P���+���G�P~ZN�7�Uv?����ϦB�Ո���ji5Ktu*g���
c�D�OEE�����jSQ��x�Ɛ�L��S��Q���@�B�}�̔��*z��ܕ����MJ��ں�����)��#����[\���.��)X�X��(Omuzv
���s�f���'���)Y��C~BB�)))�:���9��߉>>��S����kx�'�������x�95f}��\����k@C{{{�MB����i�,L���c�����D%`ߌ����l+����qJ�h��ᑫ"K ��

�@�*<dn��A���S'��l�ՠ�Qʭ�,�}⫍��b0����I�#���U���[��P��E�D�ө�pt�#��	�B>(�l����W�U�L���}<�&�g�)X���1B<�D�<u�|}��}��j��q@D�WQ��U[n�V#6��	�Eo�EO������P�~R_t�xф��2�I�7z��D�j
�;
Ld��M���S�Vm��Mu�)�����q���'5�
7\?�t�AնK-�?�,�l�Fd�Lr�~�����
LM���EI�Fj�`/~�������~�� ��?����$�D�i�N�DΜ�&���lr��9��1S:W�<����?����*��o�D����}Q=pح���mU#�s�5̄����Q6�2��ܫ��RӀ���ғ���۫����3�n3I����f��+�s@ڧ�����U6{ȿ�fFR7Ԍ@xe�##��;��fg��e�9�����F̈́ߓLk�8t.h����2�(��V�����^8�z��Y�;::�L����2�����e�jG�?s��䃆?�%+#������b��,�?�.\��V3����&�+%**�>, р�+`F�����_m�kN�m�0�����������_z|8�5F�C�G��~�7�Bc�L���+�9~���sY��/C����|�ب^��1AS��Z��-=?<�iLH�r��B���T+�ĕ<��¦'�5�"�R[�@$A;����{�DrV�==�
����7?'��x
J�s]�} pܬ� �b���~1$	D��+>Ͷ����y��5 B	~��;̥$33�����Ɏc�溛���~���ҹ%Y4Q��[�4�1��˗��z๭?sӜJg�A�H��?P}��!������Y��>Z�{�t��d�)m۰��SS��0=�����@)H����x/r+01Qii�i/:�ŀ��)y���;V��a�ʔ�.X?�z���Rf@l֚�(�V�E'V܉.H]���e`_�ӂ����u���x����T���yPR�+ �z��F/F���`�* �71�ڪ23]�=�/��ς�F����_`9�l�g�xPJ�m��{���}T/��L�捬��>��Y��000�Y�f2!�aX�`a:�4�j�� Z�
���
p�\��D1��@�Ӌ�5�T˟65�Q�'	ԝ�ڊ
�����~G	�R�o��mnlB�P��Ʈ��9u:>ڳgO��b%��K�}�%��	F��c�m�������� �o���/��y�~�q��KQ�J��D�����Ε��О��NL���D�L7�z��Y�2v���� .��O5�'��đi����g��ޱ�� S�[�t��a�{^t�9������R����Wщ�/�ݛt!򧁥�Ø�jkC-�
�������K�ɿ\�k�3 �8}�񲋇TFG��'~�4��Vy��S�D�hNNNf�/u�.p���8��������(v5Af9��s&f��� s��x�`����?mN���b�{{_���]0>g���}�ݨK���z��>�L�cߔ�|���[}��e7���'v�;�b�&�:t��9���i�w�/��$fd�����ͭ��V�קTa�|�_ex��>nb�[�U,��Cg�Sݷ��6�݁�T����NrR����20J N��������ל�n�Z*�YHgQ���)�Z]s�
�
��u��߲��~��0;?/�Z��ӡIY�@ݩ��v�{to:Yf��.��ϒ��W)���zĦ���C��#K�����
���>zt綨�|B�᫱AjUa�����{����	b�A���.8�S��'��d�I`أ��n�x"���Nxn�l�;��\'J�e�jUźM���p��*��j�>�=2>��4BE��.��KST6MJ��40H��I��LIY鮼�Nhθ�ء��..E�/rR�T�����Y�x�����b%l�!O=k�a�.����ӟ��
��+�ʳ��y�
��t������H �����q������`�
��a o�� �ȇg�G�����"�H3S���P�9TP@��%�Nd٣��+ֈ׮]�/�c��"��!QQ��<Y\LLL�����E\�1�)))]
�r�<[9�.8))�I��
����*m�,,��P�KH�)�j��9$^b��/0�F���g�_l���t{��+�+e!�&#n��N�]
���M�k}�6Ja���.$O�;��D�$�����M��Vw�uSm �[)4�C㊇2е@I6?�K:I3�C"���^�2�p�U��e_ ��g#���S5f�t��� �jX�����R[�CD2�,u����c��%v˪f�OiikgG�FQ���D){zLv�����@��&'�z:yNlLo���<�EC��Q2^<SϗQ����V~�j#y�ٺ�O|�ë�G�*�S<�ecC^]-F��y]�A�5|��7��F1�o��ݹ���6�[}ϲ�������)o��p�}���7%���}'g����R�0�����0��ü
;$'I=�M��ܭb�������lX��f��Q<}��f ����82;�~��hت��fjϴ�L�|�\HgȐ:Hľ(~�D.!�b_����rl�6I��8��}}}=111��kEe+E�:����-\Y���S�L}��NQ��\�-�H~«����\+�0�w�T듵��h8;/9\�ǥc3�f@�0j�Du�������΍5
����߀�����[�D@j��y�ر0����ݨ����U'T�P\�wx�l�p�So���a�L�ㅣ��D���I֋}°���>f��ځ�<~����a�W�ݝ2��J�^}
|���P�-=���bH[Gfi��G���[�Q�Ӌ��ߦt�����̏�E���X�,��\-=bei06�ͺ}�T�V�FU&c�]n4%���?Do�
�:�����D�ĎF����*�+üp���t�'^��L=��5H�.�������UQt����q���C��-�ȡ������4!}�ta�i�����`�6������.O|��c��@Wm�X��@�,����oy�p�]K���d��ޔ
w�9N[iߦM��g�P�9�qg5�������w�J=w	lu	����9A�ft�7um�M��45~�����48�?�(%2�"I�Dkɟ�������@;��H�;��<�?]'��I�����"��C�v�C����m�۞�mӰ���r� 	A�/K��eK�ԓK��4�R, G�/��� ���u�#�AX\HF�H�#V�f��16���]���3�/��8��t�E�MB���E4��n�XT��âj��7��A����yg��+˻[�֪�/q�ۂ���t�S�$E�+X=
��
�޼}1���jZ�ą�t��_�gzB��"`ddd���#�m֣�k/�G�ǨG�lb�Z�T�BԲ�p�䴌���oIj������f'j(���1�ݦ�d�<o̚gJB��#�����m������}L�>�a� ��T�<9�� �
�'ҳ���o/ �W�ŗ�ZXZ~�,T��f���,��ɱ���C6&��yh�^I�ux�rp��te�re(!���"���;�|�𱾾� ;���^r����*�p�v����A���["G

n_z|g�m|�;���v���ilE�Y���f1y"T��{�����IO���@����Ey�ښ뎵�z�����G(�W��^x4����D�<����c�n��!o/����y��H��ׁc|����J�t
4��uCA�醵T��v��U�<�oK��ҟ��-9e^���`�sכ�4-����d_�VC,�˞�1�XF(�2�}Y�~�ɕ�}�����7��rk��o�B��9�(�RɔS2e��P*C�$�%eJdN���<'!S��fJ�<�6{�����=��}���9������׺��p��^�c�r�OBm��P��}��e��Z[��S-mm�s̾��n�P�v��=w3��)��)A@�^-�-�e��(Jߩ#)���B����s��N��؁�Zriy9���<�5������������z��[�����oŸ�������a���P3X�}{���"�8O>z�|�2��	v�����2�W���zJ�*~`X��E'{�s�"'�Gs����b{��v&e�Qy���`?m�E��
��X&�n~A����S��W�_���H�
��{�1�8gӷ2����� ���ϳ	1�~Q{�~e�L��a�s����ŻwS��&Rw��v�Ag�*�w>����j�P?�W��r����Uor̴|���ꪆ�V<���� ��~}=�yd� �Jxǣ]�Ι���GB��j


b^��>QYڜ��id�o@J�R����_M��F���P��fG����B��4�}�t�_Q���o�Җ��9���=���.�ql�~����}!wp�|��'�5$f˸��
�]��Wz�.Q7M���W}�R���[��H��ӕ�ut����89���I�ٔ��A�<!+K䊕)wɋ��i���4��E�����z����$&�"��� BV�����ZV�G�u����ၒ��F��o���gX�/-�l:�r
���!�����݀��.�a)���rrr���m�B�yyy�^���~GڴzJX6�Ʌ]�6��{JQ�VKdXQ�d���D������^�lٗ/_���b�97����������~}{B�lc��rzz��p�������A7U����g�9�?l1���j��N���^�0A_�\Fޢ������s~%���o�g�f&>O�w��"���K��ifd����+jB縍-�d����@~i m+��o�ۻ!�_�dɮ��
��ņ��&� ���f��{�qqI8�hE�W�O7(�v�r������͒�[ШDˑN&�Df��㞎k@f�x�r��s}d���n���w��XUw�cB���{GG�_ �O-Rj��рG���*w���k����ޝģm�Uy��/^��^��&е�M*ʈ����"�j�	c{���
cH|-y2���1&f��e�����2P#j��2s*�Z��|�CB�ll2&XA=AG��pz��@U�?ۈ!��VG#Lз~7R�����v�vv���Magl:\`:,O�_pY�yzҮ��t��T:>�C��x�d�c;,uA�F&Zi��{���@<�8C;f_��J�m[2�h��j!�����ښ44
W>�?�']a/!��8�ɞ��R���o2,��K	N��P��8ٸ����	���Gl�qR���j���"�oX�>0
y��V�B�:��؇ͦ(vR}����u_��d3�U۲�/$�zn���O��H�m>ٙ�z^T�,M��� ��jnn�	I��i�٬�����-�b�)�o��[�`ڐT��M� #���:���ظ�é��A|��ɥ���餌�cc�n3���v�Ux�8�)K/h��������#*�.~rf�/z�0Vb��K���%9�<�!���E}s`��N��T�\~5f�}��>��}c/�^6 �9�ϳT�>��B�`R�GFF�I��d���0�h��mq������^��OOW���hWZB\��m�)L�����Ё�]
-	�%��ez��q`���u��
M�wY}d��>\P��X�f�*�tf�Q��I��nc�է����1�H|c�M�A�q&
RNE��ٕ������"���rc6�
P��l�oBw3/?	���!~���`͏�D�}X�1]�Y��%��
q S �s+6��Px͵�|�Fl2�파Sx�P@�XD����]fZ���YK�4NF���3��@�[�k�����*��2��M6;L��{{'���?m�"�E��.,����~YEM��>g~���.���QKH[��̝7�߽K� ����6vzD����4�a%%%�bAb��YH��9���֒�H<#>qB7�0ە8�����*�*�K��X��'?d
�LKM��E��
C �mk���p)6 ���� s~�$��a(���Ö���$�(�9i��{����n8��.R��YZJ��H�oԈ�^lo�]�.+k>��� �;Ecび�W������`cPt4G� e������Ѝ�Ǉ��4�)1L��������C���B⠖F�Z�r���>�r�p�p�7q���g�7�_\zZ9��t���s�CB/ײ9�Ǐ����R<ȯO�]�0i�}ݑ	Î���?"mw�KVN^>)�8*^�E�ig޾}�V7��q�LLL
��7o�*��6�Vn�E5��Ř`�����l9ѽ2.nX�1G���¨�ɹb��O�0�Ӄ��C��Y�b�_W�6�2�(�� �z�����#�R�'*��d��t���d�(u�`��@�zVu����s�c��cc��k6e�-����������6�S��w�HZ��aA��2-��ĩ�k�3���z�T���d�fd��#���)�ҩ�ľ>���'�����Q�v*��n���C��dX�Qf�W�2��?+�[煀���&�l5"�����Z
��A�]p�X��BэnGȨX�qd�Na�:�������ã�E�###�����	��ݻ�s���:ɐ���G��^?��͏>-��c��95]ʍS^�\c ��
h>sV5Wk���H�3N�nD7s�_, �%�az�kD��j�K� a~u0��pI��ۍ����}���^2V�3�Ȗ�(s��mN6ՉJ�����,�.*5�1ɊE66P:���$��eݰ���{�5edeA�B��>}�������p�T�QTT�%����ٙ(�������C"�sfff]��N�Ԗ�����nZ���^UX��M�AT�Qm;j!Y|�Zw����aR���!�^c����K�*?y���B�O�����UƓ'OJU��u�fV<�\iܧ����9�Wz������+D�[d�y��� B��5���1 '�d��c]<v���U>������!�E'W�)r��rF}�]f��)7�5��3�cV�AW�3`b*��a}}�I��P�uT�騨�v)��d�'���?�U����U��q^��"a�ۢ�c�z!��z*��4v;|�tV�[v�P\���,��!�0�E[C��d�y[W�`:����"�aem�~�޽ǄYb�����#�6ż�B�n���X�wd��v��^�v���x)��% ��� <DR?�<�a���wL���t��y��!�^�ƽAm��*�.
%�K�sF^V:9�'Ud���_���3�sG�V�f�g��!8J��o�I\g/���E0�N��+��A���eUU_C�փ��FZp�]E�z����!��I\�ߨv⇐(��T���ц�6[����{��m�~sGA�>˺�@^'�xs�qP7�pS���$%0q���զW\��'d��2w��n��)�Uo.��
�l��#�c�s��t�����n',$4��a]L"�׮^�l%e��q�J7;D`�h�V-�������������H�����2����/�(����p1<���c�����ˠ�O�OV���{�5��'�JouS胾�^��η��$2� �	N��q�*��i��˝�
7.���a�j��v����o�*ro��\���� ��zJ����
�444��6��~�dll�R��͂��,���x�
�yL���i�#)�����J�pUE�$߬���yyuG���z������������Xb�>qUR���qR�a�з��H;���m�A��n�t���g�;u�1gB�|��ơͳ4�J��B��}uԒf����RC0?��{�:�KdtUb�5���D��	CL��_z�7޹ߑ�nddd���Ũ��t-v����AD�r1 ��UR����z��=K e��-��;���U�? �Н;{v�ۦ::��S����e't)m�~lԦΏ�PФb���)L���D�$C���!�f�m�t?���W�a�aI���U=j��B�途��	���d��b�@��\��1X�K�0��EG[Վc�?DUs��>����OR�qJm�����^X�2�+2%;;��"���%��^fL*���XڵW��y��h����.�F$�v�v�ʕ+�l��d`�#[?q�DnxD�?����o��]��`�83�������tFw��	��a��Ν�sss#�-������RN�h)�W�lܵ���0�o��?(�ݒ�qM�$��i8Sl($p�6;�t��,������������ �~�=�7w�1�oAaa#����CNDW�ϔڎOMmp���Z��f�.]� ��בG}d��n^��0�:�+PD0y)��߸}����Q�'١��RL�H/B�:�q��@N�*����(@������I?�a�[�++�.�p���&#�x�mV�D0��5�ss��"�艜mԟ�#�=Qdە��ĹvC#'����I;���3�"�^�-J��A��/}Y��'�.�����~�ءdC=mmm3�$�1���jvJ�`ͬt���G����, ��[-
<A��Y>�����7��yR����EU�њ�5�΄'�}n�ԉ��.�X(zxT�K��}�^�����t/�mW�n���t�ꩬ���P�ރ�{���$�E���a�s���g���0��ll�\I�x��n��"��S�%�Op}Q�%?���[櫪P�b3I:!+�WY�;E�(����������+��+�Ϗ�m����6���M�6_�1���.n�]ݰ�Nڦ��|͚����K�ѫ�������S'9�	&�7YP	7�\�},�fnn�I(��(���@BO(;�!�����$!s���e�^뿏�:]x<>	�����Wr��	,�zE�m����7靖b'Kf/�V�Uoz:S�|�1lˏJ�aH܁�M�prx�(�������L4R����gT�`�Z���3�?~{��%I�8��iIɩ"�.���"hig�i�oP�4�\��A�w�j1:B029'G#҉f3 �d^�PM�\���Lۢ�,���:A�pqE��� �����@���-tD���2�Y��<EwY�rþ�.��{LF�ZQUR��{	�s��=in�a�r��#���&�ia�0��j`�=�3����<.ݹs�F�Տ�%%k`�n.�6?_��=9�]Ǳ>�f��Ԥ�4ɰ����j#N�	:�$v
�/���x�Q�y����2w�a�L5�BE{��V����Ίq�:����-��l�/G�6����)h�I;0f�2p/45��ژƽ�hg������Pj��5��k�c�`�#"БR~:ȫ�Q��T}B��FZ��d�(�FW�'UѠ�>k��c�}g	��avb}�S]�$#��_F�zH� 2��!������ٷ���/�sS�s��qֿn���3��yD@HHmYēQ:��@ڙ����EN�t"==]} �AݠǶ[G�9�ym����tO~!�D�ӧ?���a��ޠ��wu}D��o�k9^aa�"e�Y�Ѳ)A�2)���s�.Sc��޿>r��&Yu��pt��$��*�3���'$$��A\XKAA]K_N�z�9b{	ԫ[|n�C�U8�*�_���O�R�������n��{xjAn�[�7N��$j��h�KW���۠�U%ծ۲0��h���'���j�L�ݿ;2#3��W�J�)Ol{���)��}���Y�\Z�~�4��C�O��x��]�x�����Vtw� �H�c��������s�������F��]�_��F3�����\6�n��*�	�Q����� ��J������OV���l=os}�yy�8��(�̯�S���ə�T�V�a��<���������я<�m�d��o�G�Wb�=�.)=]���?��ͻ�N��:���2���~e$S����,[��Oq�d�ė/i:ڿL.��Q`��YC�I���R_B�K�6ז�>�!���5�{����샥�3{���2@��$��,l��ڄ��=K_(�0���7uiW^eI`��OI��9MB�p0mxp&z�!��}���gzT��>}+<Q���V%�4�5߂�%$$���"gƺP+�~͑�szý����K�}Wdod�U���.6���=Y���fenn�#!$���ZT����hf�$By�nԀ��h U��+�z?��x���vv{�3=b�d2� 4���#3�{���y��i.///��ں�I�g
�y>�aT�`좣���B_�����6�ކd8���vvfu_h�.EA�g�=w��c*���c��:�&���fc���-����z,�$Eg�BҞ'�#e�2�u;�8E%r�l��G�D���00� �5$4��)1�>-�	���ٳg�s�m'GI8W��G�F�p��5-Dj**�?=G�*2q		�����������.�,�6�cd>P�/��gPe��}W�/�e	�^Vv\,yh&�� �%�������n
�0�F�M�m��}v5����c2��=y�O�h\Zלh�6�/y�}���2&.���{�M�P+ŷ�6����Q�U�}�g+�c_���+�m
�D=X{|a���.S���'2C>K����Bۘ/���5�_�pQ��Q}Б`T���覈@��ӧ��I;Ĕ
�%%�$��d6��.����1�X<^�;D"��H�%LM����K׃CC}�H5!�qR���5X��v�?k3ω�N��X4>��GE���@'����܏�|�f������KNM�Dh�k�[��55���Mb_2ԉ_�h4�U�`��i��Os��4u�ŋ���������:���ä���xPż�zd���|���p��Rsuu�K��9ePp��{q�n�: t2���O!��`��'p"�˽���<�uB'MO�_"1ꡟ\�vr3g���|�h3i��������4����wf���[���,��v���_%�iU��α����	iy����;tj��>ɹ��3��%�,~ ��9$�}d=	�~��3��c�{��j]S8J[W��s48hd^�z�R�rx;�Bے����'�3Cg0LL��6sb���?�;�v��
�R�9��+P~k�l��E�@�_䖏�ξIj�?It��m������w�� ��X�[ �V�9z�9G�#�����X �?���t��`w���R�rȑed%~����X�4ڲI���{3<8��cH�����VCK��{'gh��X ��T{�c
�l�-��_Sp&#!����`V[#êf�����C�6VV����i�-mX�3������p��O�,w�w/m�{����Sss5�e��@�����W~<G�kj��'��A�fk�v�(��O��n8:6�H���YOO���%=��I�'i���~����ث���=�:�]s��ܓ	��x-���`f�@�
�ϵ����{{O@�k\��^�&����)b̓�qm���,-M�b����tP5�#8�1b��$Ύ�< -�a"�`��%&�S�\��J>DG��&=(��,���ݹ��q�f�v����y���d?
 �Ɯ_ *vv%��U���H|u�<%^t,o���'AL���BK"I�k��q-x�$��@������ƽ,Cx�@Gr���k�-[li%����,��Q1_�7�:U���\���?X�����:�ӭ7u�`�BN�/OW��+��ܜ�i%wV�MP#ik'��%pt������fR�������g�H���޼Y��e���F�퉊���B�F���ſ�E��� �i�\�k??5CK�c� �EU5ٹʌ3�d�jg��N�#���y$�JW�Ԃ��Ao�Ď��<��is�YQIɍ\;�{�ǂ0��봈'��u��+@�6G#��P�}Y{#(4��}��8=�w@_OR��ٳ��r��`���8�I^�~��%�߳4wdlL&���d��ڵlg�L�+�����5���JNS��Ps<�:_��\�O<miQ+^�Hծ��?M;)kk��C$�"Yi];<OyQN�Y�cW}^�R�8n}�G�����W�g���!��i� �@�$��m��Vؠ`���	]��J����J��h)W'Ȧ�0%�Ʒ�����	 �?"h��3�Դ��"�I0(����x��h�.����8�6�GHSM�l�ϟŃ���7��O���`*$��d���4��]��Cll�����:��w����Fx��5�����B��lY�׼}���P���㻴!T#���0�H3��`B���g^�0̮�����.;����ƍ��9�H�;�W��F��<@��1FF��'�n����ann�p:�:��w[�O⺶<Y���5��NB�.��U2:^�9'�w:�)0��6�L�/�Ҍ�V�D1���1V�^�'�yc�BRn�>1
=wί /�����h�ء��oA��]^s���Y�)oXQR��!�ͺfb�Iʉ�4OWA�!�=�FeC�
<��Ȼ-��h*6��;��S��3-�D㨣�[�c`��u@]�~|j��� <�5��=Z�vrv6�C�֑�& E@�յzB��.FZ�k�U��t����#u��	\c�+�@#�'������d���5_��>����S��}+f��G]%����v\FF�,������@nF�{C(�)��l����Vdn�X��:�`t1sh�7���Gx��.æҊ����@k�ݨ�r�q����J?|�1K�Xί4*�w(���4�s}@�BEM��p�����X�_x������`{�P寍�#+��$>Tn8��;�א8��������3R'��¨�	/�	���D��T�q�.���-]���J��7��� �s�A2bY�#�����P��㿛������'q^�6G�MԺ���ݡ?^/^�K����z�p��!;;ۧ����ʆf��mΓa8ڸ���C�w=�w砣*�([��G(ʼ�דg59ё��L-Re����e��ɧݯJ�V�	�+����6���C,�1��Y�٣�TH@/���Vz���3I�tGxA �?�_[[[��(/u���
_j4��pE������Ȑ�?����@�9�V>�ʚ��oF���r������y�����T_[ܞ�ϰ	6���a�uA"=���O*$�G��k��+��A����%�Ĭ��_ض�A��M��]汽�@0��/=�)�� 8�#rx��~�������ϥ���0��YI��[� V�w$$�.�S5l��O�Ɉq���F��t�
��<1B�f�?3Ԁ�9�od�N�gñ���!%�+�	��CO��\T��f4e�6D]k71��I���f��V�ڥa�v� �#�]�xQ ��,x��2�������Х�Ǖs��Kѩp`D������S%�W���q�Pλ���ȏŋv\���6�����doo�z�[X����D�����Qkx��>,�nr)�/�t:H����[
�9/�e�_q��g��VK����������6(�ٜ@;d���-���y�
K|A��Ȼ�{E�@pNUt`x�ЫDU��J%�Q[e�Wi8^�( >��ŋ��uoR�g$,Q?�BcF笈ܿ�=�[�t:ޭ�!i��X��#��]Fo��"�H������QQQ��,��j�^D���۷o?�O�m.t���9�}�\sI �_�|��*�>�)����$�`S���iT��گ�L�Z��'��_�"��d�"�վB|��.�-.g%����}�����Ǐ�~��:��R�1���toig���k�ܕ���P�#�J��xkm�:�tr���7�F^�*ߨU���6���N�δ�֒�Po��׭LX�`��q*ml��]��-�Ƈff�vC� ,;�~֥/s%��	B�����f iac���#�0_'{zz�moU=�6 �[��]�����FG�����r�]mNZ�d���~�����}6�`FI��ⲧ'�BM>.�c��I��V�RL�U��5idt��6Y���`����n�W t(�����/^���������_�7�:�}�����$y�ݸ<���� �WQ>�A
<�F/	���H��K;&��H��\��=��/��>�7�*�{�Z���Oo$Ε2W���N%E]*IKk��E^�{��ΝG�&;�Q6��L/��w�����A��*������zS32t�ɪ�گ�UB6�p��G\&,-*�{�$`��Lд�3"�?���������=0p�I�]O"AAAqZ\<E\N��G���6�����I�?ꖷ��>��[]]���Z��	�a����`'S�@3#3�a#:m��-�%6P��|Xe��gj�	��[�f^���"X��~�SB�0Y�E�P��9lH���2(""U\�� 3���iR���;2.���K�`���΃��Ζ��&�u���������x�s�4r��+���%Z�no�gr.��'*!
<Z��B�g�EUj��ԙ��� +}Y7�8���Ʃ
c����!���A2�q!��Z���3u�NE��p����a��s�@���4��0._�����k4���@z)Y=|���Kq�aF��vr���E3��W#�F����c�C���
������yF���]�7��%pM�>��EU��jZ��i◔���w�TlRVT��7o��Ϸ	��:�ۺ���� �0EݫW线~�ZsL-�_$��ER�K:L2B.�32����JxY����|#{q irM�{��\2`o�j�d?awd]� ȚRV6����˸bW�L�?e��Y�8�.�h�����L����1.�(����r;т<���ÇI�?#��Gg"
6ސb.��־"�d`k��TJ����H�0�Q��w�Oq��XlBm�� ��j��`)���ĎD5���r�daf�F��q���-OL�c��OMM59q��HM���^..�9�;��ˋh�H�n����b7�}�vSj�������|�|0���<`$D�|hD8���wq2�����9��3y��7,}����`�����%���QK�]*�'ܨx�����pt��v��_U:�{&�tfMCW���J0MF�n�4�:3(3;T!b�(���]7�At�.2j��~7���K2�*���v%�j�6�! ]W�X�C����nN�V[zD�㐌
4V������e�{/�����ӆ7o���Ł4�\6��a��A��j�t�;�v�43�7�e���ō��>�v[�X_��1i�z�G�ȡ��d���<K_����Z��ޙ'���3�Os=}��j}��V�3�� ��KA��Y���,�_�L%�L���ù����0��?qs�@�(S_��p���p��������*�� V�����<����gԻ��K�уebb�����|���79̫������#��19�{���֜��Y��,NV*ɢA�HoTS�H��_`���ҳ��<��������o\��j]Nڡ�ْu�Ru�j��S�����F�Y��F��$�r0,�!�<��ڙ#���ͫW9Kl2����R��$����w���PX�W�� �*���}�&�Xo��"Q'����ٙ���b�Ŕs���U2��)UM1�s����/ko����|r֋)��g���p+�O����·�Ȅ��r���������y��$�c�3,��?��T�Z�>����&`?�̞�5pKR��ІD��G�d?,^�ڵ��~oӨni|�m��m�|�=����\گ�3d&��H�#�A��$�<��8����G�>���o���-G�q{Z���{��� C�s�t{�����̟��<t�P�O�@���EU�����x�if�L�Cx���;P�>,���&��h����_�K5��{J��¿�ߗ���S:v&�w�N�B�;���.��&��:�:c����I�Â X[�$l�����b)%�n��5�ӫ��?q"���f�Œ�a��rDx���T��ڪ�"ﺳ;I%(��������޽�&uk�m����وYw���Uqϱ`%�F$#���}?/;{�@�LbtO���=l��2��΃nē�FcP���}�X�s���B���|0'V�����ƙ7ʳ6�wщTt�4m3g���/qwG�R��9�y�E�Q�T��V,r�UE>���|ff?
�n��ɗ��0%�@��sL�o\��?�b��+`,R��G��N)֓`����|:��K�����V��}Y'��ԧ����怿�y�A� n��������)��Y=��fS�#�j�ڼ�ǆ���Zߴ�}��I��k��Y��m����'9��;�.��s�[tZ�dx���(.�	[T;:#P�Yk���v>}�澞uN�ʣ����`M��S���E�<[O�������x�?KK���]�3�W���o�
-C���±���3iYd2�g�zJ�K��	X�?~�_6���?�����*c���#��a�\� ��v/�"��.T1w;=��1���,,�7�1L�L?�����sz�p���^�k6�PY���6!�������U�<�Ԉ�:��j�U�}'pddņW�q*6̹��d��2�+���Z��W`���h��jv�k\��(�Ӭ��ŰQ�#��;�NU|���2���I'���ݷOY]��,��m���zU���:���m১ꤋ��53��>����PR�,����2���t�����؃��2Ɇ�F	[�o9i>o!�V��"�x:(.�]t/�.i�s�B�^� ��I�YYW�s[�����w��?K��ܲVaS����z�"Ѫ�ȹ��t����^;�����4Ԓ'J��ӂ��`ak�N��'��)#�2�X��;�4��#�]bXp��7	?�ޒ�5��C�c�E�� (���C�`ؾ�^��>w@?�8I#��zk�IZ}CÅ��"�ݏ
3����@\��|ɁqJ����{��q�������[j�˩w�UA�^�w��R~�u��$��B���D�p�WK^!��.���`4�F�dc�E^�<�bQ��U�K"9���/��b��\��:q�gB�-:F�T�Qv��ŷ�'~�����Bx�����܇y �x���!�[�V,p���$}�R����a��j �$�H����CƆM�B�잶�]������GG�k��B�)V[}L�a�B.��Ry7�-L�R��M��z��4I�\��`�>as���x�;��T��z^�#8����A�L;�W�V�管/F�5�)�*�Tt��*(qv��/B|��dd�ON*7����1�$x�:v5#>�W���$��4��ƜxdK�}�?���h���qq�t�� [ ���ޝm�w���8���:�������	WF�ƻbx���? ݕΣ:��7�ެFItP�Y�����+�-3������n�N2"��B�o8�{zzP�y��~���ˢ�;��Ȱ?��h&\�ϟz��`�c�K�W|�U{���\�e�;�i��$�	�����	�5z�p�C�G�m��DJ,)[����{ܙ@H�ossY��Qaꡦ�~;z���s���#At�P�%>Qu}�*�:�:���/
�4��'��hϝ|�6S_l���v������5��Q����b�;���]b�\���ɢA��i���E����$ �g��B�+J�Df߆5�kE��ATWTH[$�E��g����Y��x~��N�]���\��'d��D}	Yow���A���ZM�,A��w5`f�P#<G���*�M��a\W��fC"""���4n.^�vh�.����  ((��OfŎ��&[����3��5Q���I�������ʝ�����z� ��xxV>@���1��<W�3�צƲ�H��:+���+i�1�lw���ѯ�,nό�Ta\�#�/0�WYիD͖IK4����85b>,�`����ky"�乞z�+/���x�������a�l�(��j���s�Bs���l~Os)��y����>�)�L��0ϥ��Uv8���/j�Z__<�;��`{�BI�1��o��=-"b����������O�nc�7�5��}/�^{���E����qy8��j��̖�eư"����q�fJ2D#T�",�;'{��d-r����Q���踔ޜ(>'W���1ϒ�:#&���L!�_&���j�x�OL��t���l�.���,��f�/��,K�����u��AY6�߆H\���Z^��O�8�T�*�'+-�C�)�ўp뢹���|ǎY��k��w�����F����^	����y���ջ�>ƹdHx˹����4���������]���8�ųRN�j������5����L߮r���|��G��glbbҚ���
�FZr`�A!!���֖��_���E҄��4�^�r�_;>>��!A���v9��4@R:1�?V�*��y���3��ۛE�����$Z-�z�g��W�8.U����.�lN���<>ne��'��JjG����F555�3�ӵS;&�;1c
��G43
�.�r�I������y�o���.p�ſඝ����J����et��9�eE�j���?u����;JK%N��f��<�y���"j�x��|+���SeZ�̘����5�v�h�d2����H�*@<�7�uL��7�O"L5"yq2O�Xm��1�f�к�a\E���aw�uh�Bh������_L�h���Z�Y�{�w=���W!����9:҇���^� �L0$�L�c�Lv��{hfp�_k�}a|(�e��&�ӝ����u����r���9I�v
�<L}�TT+RT�B����vK�n�������X|k�o�K��E��ܘ�y+1[�8����~�.��S����ט��X~&U��E�nuqy���J��j��{�/�щƊ��{{ �罹��>�<�ׯ����;�/��kdA(�6vo��rj!v�MP �E�j�FƐ?X�.��v�Z��gډK�tW�o�4�ZQ�U�S��ߖ/���04؃)H��ʑ:�����bO WsNZ�B7Y��qɹ*�J�LB�������������3�{��qȠS�L}þ�F)��v�j�E��Űs�IP����ϮY��x��zâ�:�?"?::���M^#��H-Rl5�{}�+V��PT������~��Ç���ϴ��I��^x��\���:Ʃ4��Li�x���~tmg�O�u��k�� ��uR��z�������.�y/<jpIB�h������r����v��P�^z�;���%Y������\\^� -��.�C6�r�6̘A�M!P���A���sSS܉82,�㶨9�{ܷ���xv�S�BR�K����+=�����=��5�<nY�.�`M���N��t󇃌Y$��(�"t�ȺDI�q�����1��nOf����3�/\踣-��s�����K��=�V=3#�'{�s
�,a��k���JU-q�/?�:�7HWL�Ƌfu����#_ć���nj�gҒ%&&~^��V���gW�w�B9w;U�8�����9�^�x���|'����4@���R'+4���4��þ���^f+:�F�ks�..f,@��t�ﾪ^�C��DJSs�ϰ�i)�����=�I�����Z+�iᱩ��~�v�cw�hAÒ��Ʉ���k��O]��v����/�c��N>˹�S%�ʉ�H�Yt9��)!G��y�I.�qn�EJ��� �z�Du��ɘ�L�[(�o��l�ۺ�6�D�DE�w�x��Q���9���i���\~&n%~�:]�T~;���Z��X�&��gwQ��� ��y06v!��T�E�N��tO�.u��6�~����軘��E��a����A�0� ��b���?�/V�$�AB�I�O/6�S{P��ӥt�^��֦&���o~�N��kO��^��>f���!��*\6�i�o�+��]?-!q��ڷ�yq����k��	ƙw��4�xJ|x�a�x�z�������qK��+����b$
j\�T���|��}#ݖ����{�d�w�ace��L��������LPp�U���̼(��@+�����񕟮�ׯ����(�	���D!���/�tF|z7�{���jJ�������]�g�5Z�lmC�{�n������o��¡�8#���Ȳ�i����JВ��b��%�7Y{�K��U:��8�����KVo&�>��ط����n�DG��&��j��#A��y��at~�;���'/���]8�?��_r�f��|a=�����������m~��4��-S_�aY��#TU�Y��xp�H�k@�AwR���Mww��K��{N<�(�	�6���ѓ��9�# ���3�Z�0J�������Z���:��Tס����ei�=J����W�n\��e���NUŗ�$�'�q_��/ �`-i�R:R��}d���i]G&7�	��>�&k&m�#�)���g3��w��(P��	q�ύ%˄�^��t-�R�duI�g_*�)w����.ǈG�O��͛7@�d)L��×��	�~~�9P���k�ܐ�ٚ��������M��W�q�*�!����y���$e#q�|qS�qZZ�my��q��2�&�deutu-llԎ����2�J�`��]�ڏ��궖�M�6�W�Ӄ9�5v��<ӟ
�@	%�.΃�q\wV�^������^��2׋s7�+�C{���z�l��� l��SF#���ˋ2�$@�띺K��O����ۅ��يtz��ң�Rx�&Z��s���>�O�}���0s���Y��bσ�Ȉ�d7�ۆf�� �����t������x���R���R��������_�ā�����XX��ef�3NĬ}Oʻ�ŢgA�nѮ5 a������3�࿷������,�P(�=��$�IdjD9C[�y�̊�&
�Hp�H��&%%]L��������I`��:���ʫ�?n�X�J�ܿ��ě&=a��Ӝ� ig677�3���;w�fDO{{��g�$����x�CCC�4�����#q�3JR�5@TA�4c+�-����XNv[�jO,h����>���g������޳t@�CZ��W����Ej_�G6��ʉ�KTJ�1N֒6�$l;Y[��է��W��\͞�%�!�C�Ǎ�~j�ظf�~/J�����~?u���_1�څ�2x�]�~�gi�`�:�X�_"_ZZZE7,y$F!di�N֊.�v���Xh<��7 kkS�j9�Z�=D����/��#~����=�7;��B\FR��^@G�
Hz�O!�m(q�z�&�2�1c�hߨ��d�����2�mz�΄ܴ ����SRr��5����I���A�,�@I\��u�$"�����<'߿���}�l�~rۯ:�d�-u�_a��;��_X�"�^|M�Q�{��qdD�Qr3>3�_�.���
��(8ʫ%��;��;����F���
^PVr����������Y��w�V�6@$�����Qf�������+����32� ��Ig�9մ���)Δǃc3����U��\���:��{������1Hk/
/��-GG�Ĥ$��:s�fl���U8-��p��s����g��u����>Rg��`��s��f%�X�<��i��9����pwe���,&Z1���Y���Ļ������G��ZwB2t��;�V�kI�k?3�3�hY~��όsh�3���}F~��+_ៀ%k���_<K��c����D팛�$g�'��2&_�ʒ�h\�u�v�l���b@���qp��.OC��w��I�b�V�͏���RK��ط��D��`i�F�WGhgd$��k�^��̇�w�__*˩��`���k5��u������;��k�IZǝy��T�O1��?�|�#��[Eϟe�g'|�οR-�@�]���j�$�]U`��u�%�0E!���{;`¹����t��'4$$��L*�u�)����P�E�F�������'2�LsK�R��1&2�K��'�5�weA�/��x��|fv[���O����&����$����N��H�1,��ΘTʿ>�1&_�[��}L�:�� ���k+D���%�ح�������ν^ԭZ+���f"A���yj���,�Sb��fKM	rL��Y +�F��~r�����c�tN�=#�D�;�p�ҡ׺��4C"�WG#����}O�/�2]���1����	��43֞�1CJ$�
�,э�;��j��Q����c<��@G���O�uRkg�_b�� �Ǥ� ������w1�`��x��艍��|��"T�� Ի�C�.X}�XçO��N�[����/���[��fEB2�H�$4�:�J���"2�d>���>��$3	I�9cI�e��%s����}��>�~�?���O{����y�Z{�T��I�eD�UceK�FYֿ0�����3���|�r�^�s'��}���Ct/�4�
R44��
O
z��9o�\�촂i���Ç��$�{q�Ƹ���
�Dv�^SW��,�/��N��I?p��	��1B?u����Ig�>�=���k]����׾��'\~��E�cg���>s/���h9�����򕔎=}4�d��x;ĥ��Ě!�)3�P��x����9(sW�=���<���.�bS��:O�����a��c��|�4(��݋Y{�v���v]y�U�r�ey��1V5Vڬц8���C졭=���7��b�/v���a���'��'X~��	.
���F& �U�R�u�a{ꭘ����)C�UG��eX
�B1�u��eN��{�a�e牚*��k�Y�������|{ ����V5�D�U��o��OY�B�:J���T��f�c��d��+���R��]�p��74�L�ܮwR�/C����$�C\��5��;�/:E91c�����%,�P�}g-�� E�层>���Q��@u�\���q�@O�`�J��b޽��_�C�WY��enm"�z�DP�ι������&�P�a��}��O���J�F���;:�v��(����70G��(��l�JY�A���	ԷIm�:&o���")ӹ���X���7 ��n��jG|?BI�t�I��f�5Ԕ+��cqc����Z}4A����~��[���<A������} v���+����N��R��M?>["��d�S��)B�ŀƽ����%�ڛ�xқA�P��n���D��!��/7p�شO�	U1��k�������7�Q���v������)|�2�D4cJ&�	r���g�'9655Mw4x\�����)U}�o��*�#Z�|�uc��3[���������P�8.�by�����6��W�=ݱI
�g�ys����N*(�b�U8@��*2x�.""l$^��(o�y\JOm�eg�-�bC�7}��,w��6�q,_G B.<C0km��M�M+��0S�s� �.��-���-t[�a����Pk�]��<�������4�=����ȇ�c��C�����v�I槁䖠�?Oi2<���~���Ʊ3g���l4I�Cg��=�I5��h��!E��СC��n��&醑�t�q��B|a�&ܧYi�Y��(��+s��B8��i���^5���{[,C�j(�Y���
P��c�sߪ"�&�x��������v�xw"Q��޸�C��$�x���"�����[_29����륕L$R�l�a�wpw���Ta �C���J�q�(�����K�!8���`qa ��7o��ҖK�����ͯp��̶O����0�a|��A �%����hCA�ER�}�gB�@}ۢD����P��ͣ�.|�4�Z)��=���e�����>�]Uyz�&�oN:��tL�ގjX>{j½[�P�>��d�!�(�_:�M y	�K��ʧF��q~��R�yGo�aB��7��|V����Yw666�ģ{���Tŀ�o>��͛n~�|�Œ�"�Ql 蘒�~,Ȁ�ĳ�C�b�|G|�V�"�ʄn��@=��G�Cf�k���0���X'a�+2�-�6{�r1��b��o��Ƕ?�<�bCb����=O��{�y����}��J�8�)5ݸẍ{�v�_���a!���&z���&�[[��?>�8�jn-Uj����㟎���V?��'t_��8tv����k���\bD��� 
�54j�2J��7(�s� �šm�ɸ�	�qy��*9,,��u�h���{۶N�����3Hg�*C+Md��(Ѡy�������ڂ�0-�0�P�$�4�z��م��Y_@@` ���8V�����L�'�E45�{.�3�{���ew`8>�f�nTm΢�B�DM�;��0���������{z(�p��ݾ}�r�S'alh��E
^u�ٹކ�~���"XxAW��G!!l��5C�ON'�v�n���;��J��tv�1Y}�cx�;J��?d���P|�ak���\�0C!��{��JU���H.�7���t�L�%�	W���c #�����Ǔ��̵P�p^�?�j�q�����o��!P�z'u�μ�t_]�=h	ЙC ��a^^T<��[����G���@
�)�e���3{���d�'s��k�J�ґg����T0t���v�Ai����h3w2W>�HZ��Ӊk���޼YrA��F�$�r#뮧E�x��xjﱁĹq<�8�̢̍��.�x=�������w0nh�#E��8@�c�/����"A|G���nx>��S���#Q��=_BB�#���TX�t߼�{�ד3�eV�s�<G�@>*�fgf
�N�am�uLsZV�M������e��;�f �o����}>Ǐ�1L]_p�����M��� ��.�wGiAk���z�t���HѦz��9�k�|��di����x�0 �;O��%�Sh�V^O�+f#�9w臩\Au����o^$��:��ޣ�f�tՙ�w	�W&�ר0��zO�߿��«��(`X)(>R�C��,�H�k	-TL�E�|�����-��L���k�9�9uNT��1���U\�
.wY�!�'��(� �P�j�m���0}+�U$���m��ܡ��t�A�HA R丝�^s=GG��>���|N{����:���=ӣ�*Z713y	q?�M���3��K�R�}�k�Y���Vf4&��h��s��x�8��˔]�<�������+�e�  +B��t�{�����B��#��\��@�$����^��i�����999%4��������F9��+զ�^Vt[���x�ڭ�����ӟ�Rꅎh"ή�k�n���$�aBL�|�7�wE/;�b-��e��9�E�k��6Y���\b����x�gs� �38�smq�'6�Oݰ�kx?�Sz�Y����wǕP���c��D0���f���)*6S�R��e4����Fu�9���J�|}AI���6 bN�i0y��I�ћT,�����_���`��	%�<���]�g�H��W�����`ff���\_����&}�H�C��� #�H]��S�#;����ݼ;xb��{��s�����������x�I�;<�	+]��k�S�i-��z���f�S���hMM���>G��Ry˯ıPƴ ��X�ęԖ��cIh�"h���`B�Z�D�è� /ZR����h;U7��/_�<8�L&�a�w�	(���7m��ц�E��_7��Tk�6��D�^应��eN��n�袜S&Vpg�~~U�6����BE���d���e=S⬾�0�Q0���'��G��ߍN�?M}���	޳�R��hK���S��)h�\�P;��*!���	j�j)��N&�t7jZ!��_�P�ᱱ\ٻ}��y�Qf�e_A��5������������Nە��#ɴ����H�qZŀ���i�=s�O�k�/��]N۝>ZS+Y.�>�-K�u��������vE2V���'~�����C�"���>I�M�3ƍ�Q �[�4O|�R����� �q)���>�O՞��r!<2r˿�.��s1U:�>�lt��a�x��}l��
�)3R��μ������t�7�9��Y��W��؇��� _"�wR1A����FʢEȖ��+!��+��#n���n��`�g	�!���ϻ��!ـ"B��d*2��Ĩ|�ɪВ{�5��ٷ�!wX���o�\==�T[[+�2�X�/�����N�B�s�DH/�FKuU�B:��"(6B-,��J��P���M���l���/(մ�M��7%��$�O�3�(a2���'��2���t�Ï���X����b%�����?�����~`��j��j��������ཝ.��e�ڒ��.� I��o�e���m�/|3u=ԉ���Rڒ���(��P�z��.Fo����/�ؠ̜���j~���8�n{���o�TRܝ��RQ	�����%
]G���n����� 2LH����O�E��o��&������O{�C/s��΁sDM�����u��c�������pd�Q-��:X㮦C�·��ь�f(���Uq ����� 5��Ҽ[d6�K8���OO�-��G7o Q}�~$��vv0���.U�u����~O'N�ٻw�&������Y����Ve,��[����yz|�ї����F�U��[̔���Z� ����en����������3�뱴9/G����t�U�	���d�oI�~�U�����99����.�-�� ��ƺ�x��m�0��0ƍ� �p�rp�4�~�gy�^+�l������$�uB�:l��!zP�h���N�qV�"[2�|��F�)�;�v����t3��5spЮ�:Ry�S�?��6��w4k����'��u�A�ީ�*��ڧ���*���+�Ų�p6�.�$QHCg�ۉE&�x��c���ƻ��~7�u]�m����7�8R
��ʃh��^]���H������P�s�NS�f*��ܥ~�?M���t(o�1���8{i��e��c2�� G�޻�Mr>�V��~�@�	
8eSc�Xh���A��g���8��ѧ�����tM�ovWKGg�0V�[H�ZD��,r���__��I}�q(���=f�A�?/,�vP�G��,�T��)�9��h��Ŏ������[���l�r���p�hL}>���I����E���v(iW���B�>eɾ��Ln���>z������(��˹Of,������/�[x��|8�*��2���?�p�2L�ծ|���Mh����7>����I^�]j�~,��E|��^���D��$��L�D��z�š��T�@��nS����ꮵL*?:FB<���v/Ї�F�5�<*h6GE<{&����g�`�%����.�;�[��H�2��:D�h���E�Xp�U�Ĕ��M����vS����A�?�����8�`��V,�֔�^@�
����L�ӧ��`�m(_��-M�5"	�A�i����Lè6;��r{onffV��Z�?��?��ն ��ZrS���&]
��t��2�y䪁��,8�8~:,N4������?w�]�r劁���4����@��

�  ;�����Q�^����cV�,�
������3_�E��-h���c�/�=�JQ���	3|��H�&��3�HO���(���x������.����W���
p��t�c��b�K��	����6�:a��}�Uߧ���M��3�L�&�N؁4@8V�AB���`��?{Ai���NXUc����?E�I���"�����5�OgӔ�E�-��b�ʣބ�kDR�W�Пb���uz*�#����o^rO����aɲ��a�E�MI��$��ڝ��J�}r2
N���đ#>J1mJ����y�+�v������R����D-E�h�|�Z�5]��^*A��:4�}�7=da��hv �{o��v��[G��l�sҗk8c�C�b�s�S�ۗ?� �	Qjv�l����7T�0Q(Fʾ2�P���w�&y�����\I�H�A�O�0.�����s��m#*Q\��&ܾf9�A\��c�m8���	P�1�Q]�[�{y�c �]2h�o߼9��c�P�� W�����ׯKt3�v�>��Șxt|��.�6��󫺜�^Χ�߮�e����rX↫�bό�܎ߕ������g`Ԛ�g/���S�/��>��M�thF�ǟ��.K�(;,
��#9�tV��|Z
#��-c*���]!݇��ų^;�ݻ+X�b��~J~c���3(��P',�;:A-4N#�@B��"s����5�gh�d?d����K�K�=��b�|�����x��G�0M�6�(em-b�L��i���"U�S���M�V���&	;�]-��(��)��9)�� �`�yl��v�kt���}J���p���6��Ս5ճK�O[�O��[�S!��t��44�:�s��Ѻs���>����MMg��}� ��ψ��^�#`�1����|�@oZ�o�Ώ�2���w��{Χ�xo���Im1LoMQ�����̥4���Fb�P�WZ<9��[�a��s�4�&�Ɨ��1)L�>5�&�C�]�Ɵ]A��[+����P��n�7�o���8������)s��'k�h*��6JJyb����g���}�k����I�^i���楛��Q�s�Jqb6o�*��-�A(��r�8V(�X��s(=�N���XIa�k�ǽ%�T3�׾�é�����O �|�M�;���ף	Y��_!P��E]7���O/�$�+Ҋ����J�[;�O�	d�^��Y���1x�q\|��^�.�ݎ=W�Z]���z�F��\��:]�}M���]a���V�)� ۮOd���^��|#�����?���%�L;&,HM9l��>U0/��E	�+���b���o:^L��⤟�ʧ��Ģ6#O���D�$����;�/�T��rB,��arӗ �����}�-��^�	P��%F,}7#�oAv[4�}�|���0@I=@J����s��s�t��b���5eĿ9{pҟ����4|���Sn\Zz0%#[�'�E��1%��h>H��T�����ع�y��tWee偃P�n�]$�qHg.��z�=��*���i�u�����هJ �H�P�.�p��gƬ������@-RFJh�<����_C)�pu���K}���M�~ʺHf���z��9߅J�����W��Pc����bn������!��L➔�$x�g���rl�׾ۭ���4f�=?�o��Yve�r�xO��Z���z�Bb���@�����a�<<<&j4X� >�7��;��R����� u�in,�&i�[CO��11=&��l�6SNb.v����@�+�L5�X�v����;6�`^Hƀ��Z$b��V:g�wRfo�L"�~�Yn��{��C9)����f��k��Y��;��s���Sv�*B��b#Q75]\��{:6�l����up�x���� �/���?�U\�S[H��(��,�H�� �"��{����g]u�ul���V������W����������(P9#,c�J<(�e��1��&𢳂����NY���`�������|�֯߸q#�Ѷ+���}FLI3-#���N��$/�F�B?��KJ_4����Ha�9�3�1�,�`��D�;s�B��$�[���;P��j��������~(�����C @P:=����1�/�qc`���rUW�Lހ��B�yf��[�j���\������/^��A�d�";�-k�m�GSr�����G��O`�{�U�?����SH�O+:@Á��E4���.���g
:'�oE��\[��J��	��-[����X!�L�O��B�Rcu�ӕ��Itx��`'z������� ����������
&Y8�ńu<==��SF�MPO6(��0���
9����,z��3�O2��S�
�oҌ��X���U� Q}}�� ���|� �V!�CK�a9��h��)40 ��޽{��{��5�#�B~`̫��k�aAV��O��u�/�8Td�8�3:�	��2����K2;�>TW��=��,�RĲ �l��u��Kn?���ˇ�4\����>t�ڶ1oӸ��Q�{��_�A����D�4^x��6}j�
�X�������+��:b�rE�7� 1i���8`�/ۧ�ԏ�]*L�ͧ����>��b��1%j�����e�bt�~\�l�{,MM,YIh��1F%q0�_oH$1���x�$���?�;Z��tu�v��䁻����Ǆ[k*X�u�N\1�a�w9���ݟN��(~�ʛ'6h5Sį��S���I��7��� [ <V��m�h�#�K�:՝�{ک()t�3~i��R�����A��'^AY:²i�җ�#�
^��6��C�ס�5��ƫ�Ԋ{��):�>��ϔ�p�����:��7`�����g蟧7���p��G�;�Y�w��K<4EG_�AO��4o��Qz�@|�>Ȩ�jFFFÒk�$/�i�LW
�efh�v�
�����g��<�P}�v�W����P7ύA:E}�357l��ɷ�?iI��81cJ��gg������M��XW�J��X�����Í���>a��Q�'C�f:�/=ٹb��:##U��ö��,Qa5��4J�>II�錬���O���J� 㜅95&� 0b�EF�↟7��n�v�K-�bjU�q�⩅_վ�ƽ�6�&�nH�|��H���g�F���Æ�̝���İ�`0�G�w�����_�g�IiMⅪ��WԂ��:��3tR/ ���&�DlS��ˇ���m��j�,�e���soR� hu����ཿ�Zgz�>s�t����e;��v��Y�5�OS��׈U�"sv��J�؟M����@t4�7�ܹ�x��<#5<�׈�M�'_�t�{.�q5���!�/�͹��(�b+��{�^3��Ore�l���A�:	r9�j)���>�R�@8�(�Ռ�~�ج�;�MEE�?��B�c�n��@h*,�ȳjK/����k �}�����U����ڄ�%�7^�J��K=P;���j��̲�Ϩ��^�}�2a#F��xr]�o�Պ�ske�*�"¯W<o=����zZ�g?:g�O����|�q[9��N�hoݼ�v�t�"tÕi���C�x������3x.����X9)��1�i7,�;���*�j!eܐ��Łv0G> �u^=O�vʴ�'P��r(���|�+�l:��G��[�V��i0���6(��aJn�\���\��(*��*������k�����l�ɻO�����\i�Eі�t?I9�a����T3Wa��T���02U�R5(.Q1y �֓L/�G!cm�	��r(�R�aoG����:�<���]�R���5�٪ڻ/�p��}7�8�ܛ!�	������)��[	�6��m��
��a��sV:��ь��u='E�x���j�-? ���1qQ�'�����y���g�	��E�Tt���������PV/������$���Kܷ�/8��鷛�@b�g�ەM��.YkI9*/��0�ӕ�h��aۑ�嵳B�3gX6/��1�d=�U�'�!�K�]+�fjcsv��`����E���1.��B�P�Iy|CT-�)Y3�l����)}W�s�'�lz�W���'��=;��NȺ�}���S���v�s��ϖY�X5�&D��ާ��F�u*m���\���1m��Ͳ5�RV�K�cs�{Δ�f���V>�kݳ���S�k!�Fv�\6��\�yA(��{�����H(��ϟ?��ҫ+�=��z�J��nV�
�"���r��QUZ�iU?&'�=�Kq����N�R�dpPP�-�߆l�A3��:�{��Jl�	TDy��ɽ��$�;#B�߳ ��RQ����w�f?�t�P�DM�3�y+�}�������**TJ�o��ޟW��S�� ����"�pCğ���xw!�F�oe��W={�,;���$3&�{��\���ccc{�5����.꒺���,]9�Ӱ�b��[H���,.\4�q��W�d�����y�ܡm�6]��$4��';���@���o޼�0��+:��5h�{�Х���OHB9�R�8���Nd�_�q�(�q��EAy�L�ԭȶ�<�Z���_c�ϴD���"�Z�u떰z�[�����W�9�8؞����C,�<�rߋ@����M_W�QLN��JI���jȐ3 }Сqѻ&�����a� ׅ�~^�J�Z���y5�#L�De4�w��t��~"�%<3.E/��El��)L�̷�P����"�}nhh�e������J���A|��&ܞ/P�'U���r�`���Yo�VDo����P�Âo�rrr
����v�t�X-�s�C~����s��F�8��#��)���`aaQP�t��e���(�x*Q�:�@O��p�%S�� �s_�b�����v}��ou#�oIW�3%��7�?���t.�	x�PTt�L�u2�pin�d��ܤ@y`X�4�j�	���A�4��{��D�U0�"Y�EE��.��D����0�De����/�9zk�QSe�U�۫���C:c2�/�L?~ܹ��z$h'̂@�r��M�TO��ZW�OB����AZ��wIg#�f����N����EN!�����H@�3(�ܴ����� 1�PNU��	+��X��l�5���~���p�S���&h�}z픪��=Ff�e�՚����\��v\!�G=m�|~�!yHv;� ���gE
j $^�WU�\3a�^�E(�r��1��-��gI�*�Hm�����8{І[��>����]'�Ji�j]T�����m�҈
@�NC�A8�pl���jjj*���t���}M�/�Z��f�$�����&Q�(+~�����ڵ!{v�u�E�?h 6Pj$����kޠx��"ڪOi~�V�ld�Z�3�۷#�Pc�|af�ۃk�m�?���c����ģe�B ��������X���;?�!��Ec�� �#�ǅ2l�;�TXݻUUU�GB���+,2`qI����>ǥ�CO�rba{96��y����/[|�6��t��Uy!����ˈ�)){�h+Z�	o�e�Z�!��V��/��.�@��	c%211�v�?KJ���񹦇jH�H����Gb��<�C�~^Z*-��R��Xd`>VbL�}]���c�q�Ͽ�tz7A�u���\�^�:?B�����țe�v�X��w[M�1�8gu��=O9�\�.#&q�Ȩ�3��jdaj 5�z��F=��D�]4Rt����*�L.���v�.��"HV1^]���Ʌ�Z�t�::�ҴD��~6���*x���+����Wv�7
���J��׳Gh��f ���5Q�h!*Ѽ�D�����l�{����@[� Ꚛ���۾Qa�2��F9��d��q&��	HGq';�����NEA!^|�V�LM��zIÏ#����"�%늯է�:�<ڽ��Ô����Z~m�Ny@A�~�?���햣㕲��GN|�����B�a2��)�|S��]X�t���z����w�i��s��k�츹���O?���VK��e�_%�m��S���V�i�K3��HVj�J ��I�T�GTJ��\����p��ql��;/k��~�\�¼.�~�0!�m=�4޽G5x;:�c��r�wŃή�������!�����@�����h`i:b"؅�c�y��{�rrr<�G�m�:-0��^�p'�v
Z{ �*�1Լ=,�2I��6(/��ý�,��+�i����2�~�v������G��������q�-W��._�I*^�PM��я?dƐ��=���C��T�ڰJ��Ȥ�BU��z �q� $z���gUDr455oւth5��0�W�\Y(�"�H�3@�5a��Pf.;!����(W�B�Y��A�]0��w։?\8,/���ݻ�;���R��fׯ�H�:0��J����{p�0�\^�����	Nl�ɒ������j�����8�_fA)��2}ii	mhM&����/3�{����T�!W`�\`�����e�8���c'��� O����K	�Jx�y,6dBzXe��{������ێV�&�@�= ���n�ӧO�'NT:�;_�4@�T�
^����������߫�*j������7QVA�Y�:��YRG*B�t���Ѧ:&�B�r�i���߉�|9h@-E�k=���A��qqj|��$9�7�N�$2��u:Q;�^E�-''�,�e|��By��0K?�'LW���s]��t@p5���(�.�)*^�h}�a���?�HށR���_�v&��!SQs(	�"�4\���ϣ1T��܅	?W�}��������<�f��K�O�dd�-.�¤5�VĿ���r��C���J��}BQ�����i�ɦ��e��(��bP�.)y�4�L�.�h����,rw%*�̆�~��GC��C���.�������Ֆ>���
���Ʉ��++k?�O�Y�J�P��+Lf�i7���/<<<�V�X�@��(E`e��է�u���n;�إ,�OȢھ7e-6�oh����1fʃ�5�ep#y,�8?����ߔ�r�$Y�k�j`����-�*�#"#O<�vŎ[��W(d������'� ����)	�@ �������T��,DNg��+�m���������){��Մ."0[8s�Ν�Cu�G�䅲Oo@�V2@$��t�:�k]���4&E����rl�y��P0��B{�8�Q�>��??��x��R!��a��/�n�by(����F;�b@�R�
<;�&
Kj�T/y(w���X��;�������E����7フ�����}\p���.F��.�6~D���-�T�E7��%}J�B�����<�NO4`}0z3(�smسW�@���G�}r�m�d5�FVQQ-�fJ�WI C�l��<xH�Y]��1rG
�mT�����Ż�:H�+�F��444��<<E��u�^C��H�bZ��5�����ܠԒu�v�=��$�%rC[�s��dL:˪M��`�ړ��k�P#w�:�y5b��6xʅ��L:{�;oJ�9ev�g��Z����F����p�\��-��87�Jn��}�����#��'Z|YGG��xJ~���p�d"�o��s"�n�Ӌ����_����kmC�7$1qWxLL+%��[��쨔�E�4��8�g54������V�YX�"�aԻ�kZF��:��9�~��Q+Y^bq�V�����������N��4e!d��!��烂
����h�����U�����j�X���"�;d՛�D�Okj�ˢ=-�~$��O0��FF}eYYY��EV�k�"���=v?6���^�3�_�� A���ߙ\�"	L�6��W�g`�ָ"�����9Y�n��s8z��
�В����K�s�rσ������wƮ�2O]�����;;eK���y�a�t6���!���ώ�
#�-�㲍~�l�B�f��|�ف���i����5?GG�V��s*|�UY]ɶܾ0�=���B�>�Θ�i�S,�U�^M���=����w���U�KAU3��`�����������
���_��I�&tƐ?S�>rS�k�qFo��h,�8��u$��d��V\�x��4��\���J��9���Ĉr����D]o��c\��.�(�)c��u���~+���'�t��h��}Q5b�����Mm��r��B�)�(�%�--�����i1N�=@�����g�/��o4�t�q�뺹�����|�1�\���~���0��e������'('J����(i]Ӛ��:�Ef9�-~�����>�<V1F��
�v�� o���쬼������.���2b�8jel�T#��װFdU��e1�p���ؿtpv	���o	]��)�| ���7����z�d`����=�v���ȺN��)�OH8W6i*����j


jcW>Ţ����#	�zU�S���V�r�$�%�7��:�{q�S�"��s�z�_�L�[�,7���1���0���Ȧ�W��Aló�Vm��V�9ڕ� m����K	���]�}�荏2� eT,�5��[��ъs�W�&$$$9�ϻv�'�F_�i~=2(N
�2�!<c <c����68h�"�|ӛЍ�b��JF^�s���z��鱦�bRYY�;�����%��F���*�a��؂��*�&��qv��t+��u/�o�5�zH�V�c��H���c�Y&�*�ݗ���/��,tNO;�!f�
��c(�����9��ܗ�&<�����;�̓DN�u�SJH��
�c�9�M��������o��#Se���B�FZw#q��:�����*[���u��ա:���Ű��6^�ԕ}mr�?}�ܬ�����5�z	���M�_%��L��:r��Q�m=����>��w�ЍLu�+�*l��s�O.�m/(__�����+�/��vtv���m��jk�j���V&�a�)tf��̕+�N�2W9�j"4�T�
��,�u�;_��x�r��@�ce]�u��'3��߿�:
Dk@uDVi��7�~�e�����a�"��o�CC���5�@f%����$�*İ`�M���g��G~�0����5!Ѝm���쏼巽��
�R��Z�u�I_n�|׹��nu�#�|�m����9DgF�{�J��-� �THg�#�>�^�q� �u�	֮,]k]$������f 1��[�Q\��\!�vAL��"�@����e�D9��A�H{�L�	�����������`�96nB|��W���v���ߵB��IѾD�څ��C22��h��?X�9a��a۷����://�h��7�[F:����Ѽݶ�������^�z�!�bq_]]]|PP��k9~�v�+Ê����QN�d�v�V��BUb������b>�n���r�H���и�g [�EE�^��2��T_��;�҉e��Zt֐t��ҏ�к늑�Mh۰	�RJǭ���j}�e�I4�t7��17}�r�9� 6*,ni��ݯ���<��1������@�^cy��	Wz;;�:z{{��}Ky��>,T]aᓭF�Z7�ˋ
�77���j�wdV a��j$bw_w�t�/�.(�S�|���^ƹȍ�,T+*$�R:r���w%�5��s�o߾�B'2k�89ss�l[�l���'������h9(��'��N-D8Pj�&�{�3�o�:Vdۮ��ǿ������N�M��L�X���9��-߸�]ЫHs1lw��������7w D�s�n�j�~<+@)$ꊃ�J��)��G�j��w�޹,'!9y8�M��TdWA���~�>����;����/��DQ�u-��*�U�����������������9yC*��<ȃ+)�)�����w%O/�T�,�ބx��iXX^��1?�G  �� ���Ǉ.��3����2^�Ҏm���c$M?�V,`�i�%sJ��{?#&&�0�oA,��y�ЈhD-ܲ���F���"�+��P�d�g�C��Ô8�@��1�'R��_�j�J7Yzx������i�4|��-,-m� �O����*����GgTL�s��Ҍ>����q���<LI�O>��
�/�3��B����z��37�:#S:����s5�&3�o��Wx�ܙ��p��:���~"�s�˓�z�fn��?.N�V���]�J��Ĵ-�
�%2����8 �
Ed_�
� �mba�]C�^�5��[��=���mX��t�� 6��Xmړ�|O����>t�<�j�@�.��VVJ��www�ڎ�ؔt6�u�zxD�W㚁�B��@N����ݤY�7��C&�!Y�se*)$�-�{�7��ܜڴ��PX-�g�|�}䟛p��Fzȵ��J�[@��9~$o�A���ѧ�l4�;0Ì������W{zz&V:��8�l�	Lۿ��~�5Q���wܼy��תZ.&�+��54�x¢��@��6���ޑ��d�Igz@������d�:��08��5?�U�
��r"WP���}E	���ryw0&[��!��2{jj��vR��'ܾ;�P���
A&�D l�f�s��`���4��2oZ[��{��3tK5�g�WvGp	��B��|«��Z���O�m1P�/�D��$[Klu�S�����w��DF!�@�����`Z�F��w&�u|ij�Q����+�[��Kp�hy�Ɍ)$�?��{쑚0�E��Z�>\[A���o�q6�;���H�q*Qfl�.5⤤
�?}�|��.���"�q_I���M�![�[[wo��$��h��D4̻�$��D�{o�E+�fw��IpNֽ%EB�0OëzOW�����b��l���Tm�"�HMM��ⵕ�u�х�K=q��o�fgg�K�e!,B��n
h� �>������I�&}<�n�����,/��w�Uzْ%`ػS��L�*Ӭ+Ũ]з�Z�\YC̑���n�Ik��}��.� �§�a�����6C�/�2��	��1�O��?��b�KZG
a�`�`̙������"""�S�#�?�O�����l� 6l�6d$aec�zK&����|�39��9qμ��V��Pp)e=P���ܸ�J�w�	.[&Pa�<��+˺+��*U�)�-�{��@�ʷ@��1l2D��Z�r7OO���E�� d�:PW�3����f���]?$!Z;Dه���a�r�,p�M�ʮ�Ȑl�������{m����H�#O&��c��~�h��:�3QZ`���l�����t�����fRp���G~w:�=R����(��̕u�w"�Y���x2@Yh��v�	�~y;��;��n�4��@[�i��ߦ
!M�_�'���5+Hٌ��� bFw���p�rQ� � m ��(�7^�fXc�k(o�M��m[ս/L� 6�	dKs����u+`�Һ�=�U����Y��������fff:��Z��ml����逜��y
����N��g����ٳ�����<�]���&?0�<>��d���F4�:��P�m��	�pX��/�z��B7��5�����63�LIMm����ĉT����j��������ͷ9#���#�9O�}���`Z1�c���|}�������B+ƌ֗�v��s�,�Ց��8z�Rjvv3Q�����8�	) ˫ff/L�/��rV�|��uGv�sO.�b�>V�S���yB�Ω����"�1+M�t��I�KJZ�S��O������Ņn2 "}�E�bPf�R���~��������<�_��Y��/�� ��Ξ�(��M�ɏ�/!��2??;�.Y��8��l�/ 0���H�W�zT��OF���#����M��)� K\~��I�������0��:e�XR�-nac���4�3MNLAE��V��\�^�#V۳
�:q��N�=ߘxŖ�����6���X�ʜ�������)�n�Iq�_�R�C�m�,�@;�;w�,�
��،�57�����@:�����~P�+�7+*��B��������a���ͦႎ���`/����	�#��\����Ω�`X���I���~m6.@Z k��A��şaaa���e��{�Q����n��v����GDV���,A)|�5�ci���G�P�C���'&��nnu����'��Y.������0F�[_���u�վ3Y#z�}�l�k�D�W ��ܗ�w���Pځ�1US�#�����E�iik;���`��ѻ����g��l���Ot(?�k�Ov�&pˊ��4�����GGG�'4%�M-W�`n��%A]��fV����JO��y�?�6�`/��΢0Zo��G����^i��b,��zOKK��cQ��t�l�>TBw(R���U����^���VDa*�	=%���'�8��,�L�j��㟃���0(���jN?��� ~�䂡kV�H�M�8L��n}sX�ӯg(|�c>�5�8�|^��СC���<V����B�����:���eä�%�}e����_x
i� �^F����+�&�H�xې,Dyм�,���]�[��+M�j-�<��Rg�����J��}=���{,5��wY�a��5�ͅ�&/��2m�0C �fw���R(���M(k-�%�Y��	X�;Ӄ�z4����Xjc[���� 8�8	�*--E!���uL��(#:Ћ����9�o|�H����������W�&���ݷw{�+,��PpZ�ь�Ҝ �L�u�������f>U(��Kq��?e�Rذ��K�sw�@�Z](6�ˁB��8�D�m�^8&���\���"`��K]�}
���"j���"�#������Pk�E0%%�9�:�dP{�!��
*j��3�60&�ZM(�*�-�����t���h���=���g��ɠ˾�������뫷�ym�%Q�
����/���kk+�@�<t� �F$!�:��Qõ���}vUM�=�N�-�|@��=�.����eSA��}�w�7<>�n�ӸAĤ� "`]���$p�in��J�+R�'@8��Ԁ�i���$j�be�*w�i�Ang����{�.>n����apۮk��}��ڳT�]{��Ɩ�@xl����]�q����t��#J���4{z�Τ�"��~G%�#!��QQO(f���i��[!%UJ���t�-��?jz.5흟�[O�����+u_����Kd��M����ýͺ�U�Ut��%O�����0��� �ƲA;++Q�tNZ�>�}�m������DP����33�J�4JR��n	{����765�8��{�N���=7+l쯄ErG������6�O�M8@�8!^�oi�t2���8p�]�Wx��*���\d@���/��N{w@�{N��rozz:R� �G''�.����տ��TSw�mAc�m?��9���/l���~"��'3m�Jr#�Ig�n��We�s�O����MLNF�0��!j�7c����s���111���4ea��ZOM>B�d�e�S��`��P����\���4d�'Ǽ!}t~�H�a��}� �+�$��䬡�V���a���]QU|�j�5��-�,?��B����б�Q�M\�`���ǉ> �H6�t�y<W��?~�ceȐ2�(	E#�UIҤR�\D��Ǘ���J�����<�%�Jɬ�)������{����w��✳�^빞ϵ�^7Gjj2�암/x�L��)`�њP�ì� JaB��7�-Xº���-�7oƊ����d �D6䭂���9�n��Ė͍�tg���h��&F8�j�֟Q�������/��p�͛�2���J�/���{��t'����o�%��c�h�������M<P�y�d!���r�ʧݫ9/�8W��Ǧ>��.���e����XL��-����~�MoCP&Kr��:�㾞��p������r�E�"2l����TbN1'$]M���2�������t�X�>||UY�ܷ7��0�+O'�����3Q'srr�����ZZ�������8.y�έ[ �6u�M�&x^"�lĮ��l��/���L�`��n�0Lz���A�M2Sϳ�8|3�қ7o�q(A����^̼��{r=m���Y�u<�>})t�,=�z/���w��:+��ח!��5O�}���b��cM�쟷�a:�2xUx���ԣ�/�3K3[�(��4�_���p��;Sl4Jdn`�s]��N��82�y�!̢) ����N��J``�'5��!!/LX{>���707�3+f��c�/�����+4�<\]�����*�:�9$�FF�HO�G�0]k���ב� W�Hy��{��-:*
��z,��Ȝ'�{�W�n;�9���`ooc���Ec�^��,X�hJ<2�tyd�WPa30�3�Kh��5
k�������r������j��������y�mJ�l�1
�WQx񻳄�~�����d���>�ۧ3����Z�d&�`񝟳�;M�֟�\f�����y�������R���bf�L���+wDD�S�ut�t��ݻ/gvض��̧���F wǕ�:��w��gW������X�����bz&�x����$ ��5�9���V�����^Jf�J�޽�v^���b�Ǎ�%o�p�8l�>s����wtT\�{ ^�y�g�+?4,����E��5�Q�Q��S�Þ�T�a V��1�@�_֫��֛y�5��1��FQ�q�^��	ZR��S��?���;J�[��orQ��*L�l~���[���X3��N:�+"�� RN��'A5�^��`�}��L���Zu}�^]��z�x�Yb(ÞݟʾY�sY�$�aV�����^b�v��tN����f�"Z �SR�l�N�Am�h٧��6ܭ��edhxMK�������D�FYﲱIO�3ѐpCz��?��Ƅ㳠m���l��Z�6 
�ь�����`n�G�`��X�x��AF���S�ab�{�b��Q/4�_�B"�Բ2��L�����C�ǻt0˩_�ӓ�g�[pz����yc��||JE��X�p
�3�$n���_Kd��_�k*Yt!����Ա��!���.��.@%�K:��w�N��j����m(�ɓ���Į�5�y���b�m�����#Nɡm��Z��C�v_�>z"�2���`��1�2�~���h+ƪ3g������ Z�O�ޅ��i��.�eXr@k�;�nK�[Z.5{i��J��'0{zzb]�hÆG�\��v��"}B��纫~W�����}`H����c��)���J�Uvz߼�3��f�x]}������Z�e��~S����m�j3����Gi�(9���uߧ���fY���*�1-�i���sÕ�U�m��~�Ճ���1���O.p��b���K��T	�B��I�u?_l)꽏)�l��0΀���̏}pp^Brjꮧ_T$9�9o8lhNj!�ߦe�yX[w�HgW��n��iĽ�m0
��G&��7������K��ȼ�aPF�R���:�k��R̈jI���M@,Nxf	��|&��ݥ���TM�vuu)|$<�y���L؈8����z�L�s堙�qfFF�������:�'�����(�� ��1���@�f5�v�<�sb�1�@W�mw��;��%ݴx�2^_�ښ%+��.eq�$�)����K��C{��n��:���鉔i�쬣5��͕q#	���L��Or�3���}�G��;?��z�CA�T��o(	\'�j�
Кx"��5�8�������R�n���0P��`�5�����c#�����˰�q@8�?�{X���&�_)����?���Vll!fY (Eur��$xF�GY�,��*�<ZVMyv�ud�� x��ao�[�56��:<�/}�w�f^XG�x깾�����tl9�y31�x��ΰW��m$7_�ИD�m����a�����Ǻj��G}qkno��ѯ4��K��uu������c�>HKK[��,q�Q�ܨ�vrIŮ����[�T�鮹u��p#��P���&�~?�p�zo��M����"��+� ]lה6#<����і����&+P	r��P����۽�d�7T�Jg�z��z>�c�^��M�'A���0��z�;U��"�s:�17���}}/����y�\P�������.��0��=�"�Q���rڪ5���?hcc㓪_�W�}�l�;�%�7���:����)53s�ˊ�$�x^m}366���|���{��6�_����Fa��W�=$̚���<io�bq�h��k���'>)
�T
U5��R�����-�}q[�#��$����=��_��,"�T�#�d�{8oq��'Ņ� "�^h���Z"=q*41�R^P`�$@��6��� ��7ΣbM�|��b��מ���}�L=��q�+����<�&����T��)N�NΗс1;�W�	JӠ�����IPi��#ǚ~?h���o�L\\r�CO/�B'�zu<���8\z�dk߆j	�������N!%����u��!����+�Vf����EdFs9�r�N����8�k@���O�ٖ��6���N:��3q8��Y`�i�\!��q��Z%4��=��j�27�;����͛��v��h���.��Z�3>@���J׬,�YtU�:X;�K�a�顱5���K��ZO����.H|���la�0Xʙ&Ԅ���	��;(I�����'��^�Da&`�L�oS��,��t����*���b��"��Y�g�3=���P�"�_}z�dȫ��{�f9vh���|,Hzӭ=��C[��E�6�h��LX�MK��c�(�E�5Hi&��g��L0��vM�R��~\���e�ec/�,�>���B�O����O���U��ڦ$}�W�n��������I��Gx�K�y�u�=~�sة���>�f9u�Þߤ����6}��1#�#ʫV�b��`d�KM�c5A}��,9wq�yX�M�k�z��xl�[�1<~�Ҕ�V_�W��O�@dh#�:?��wЖ-�f��rj\D�����<���K��:�t׀���@v����5v����i@9R+��dr�:t(��&]Xr%�+Nj�
�C_���>�,#텍�5����Ɣ�N�ev���&o;��7т�Gse�;X�7E	x�4�Y.:x���
z�MMLҏq%Ԑ�'�'=<�\se)yQ�L_�EN�{�lI��H�`����g�}�t���2W�������v�\3R*��UO{�a����ǲ���t^�R"����m�#�dX������l�ו"u�B�We�����ʈ�f;hlK�_�e�wR�-����~�x����L��h��`޷o�Qȹ2޺}~�ׇ�V������#ēP��<͞��ќ�8*3z`��^�؍p�汝1`[v@#]��������;�&���h��ܔ˺��x���'0?1XR������&����z`��911�������q��;�_>���/4�of9ٚ�w������q�N`Y8���t�\ ��%��ݾ�Ed� ��rT��l�_�`3?k��e����%��.a��!�k:���V�:��%�-���iSM��10<�F�<���Vq^#��Lz�5 :���ug>�0:/�����ɑ�2��ϖ���<�������0p��K�]����8���A�k����@�ͳ�^c�}ڦg���ݷ�_���o�����r�Œ�Q�O�Ftg�:���v}�)6�:e$�Q�?�V)����+[GG�A;��e��/�͡�������b��]�m�>���<��D}� r��q��7�~M���[�a�<],.�M6Q�j�/�ê���5W!@�V��q<� |}ު���̄ԫ�]٘73�/�7��x�>�&�SI`�4;nvz}������DUue��:�66����/O��*b~	�?�h��R��M�;��I���J������JC����0i�W �(����眼/(Wsg82��ҋcA����:Ty0��ڪ�2S��r���M�@8��Ivo�l�$_�y��gU7nL�%X糸�8}:�0*)v�UA�|}755%�W�=='�g������&|�:�f	
�m�g)��e�"��DY�	�?L:�݈?x�L�G�ihu��X_|�򥕇��4��00uۅ����4 b8C��b��3�Y>>Q������u� �-HC>�h%��i���b˺㏷�����"��6�4�r(�H�����l�k�����8""�-[qeZK@��~`�3ہC0?4T|r�+59�=�s�=5� 4(V|~恥��}F����z7�ȋ%�bi��f��-@I-������������O������rHT��tTDXX���s$���]){c�A$�x�by���}@~n]����ǘ��6@�u��%ެ�P�h�_�ŉ��&x][��s��yV�~�涸�^҂��5��g��/��JQ�D(����J�f	�H�/�Yb���g
b�3߆����|�I�|�S����:��� ����� �?�?77����3�^�{F�������,gΜy�e�fmd���I����ێ�������~h��<S!��J��T|���NCوJڂ�Z�q�غk4��sx�ǯ�і�Ee媟?������?<����M�Ӕ(�aG�s���?����:�a�����6��b�g�F`u�H�l%W���� 6LS���mj^c._�J�l{��tfx�>����`�-�ӇƖ�\Z���&{`��P�VX1w�`���\��7<���ӷ��iS���>m��ŵぁ����� ��á	k�"���=�{�+���������@��odp���Y99��ѫ��s��@��P �k���h��srrr�F�������M���oP�X�a�h#���s��߇;o��h�_Ϋ?}p� ��-��T{x 
�[�ח �׹����=YvDF�E��i����Vt^���W+o�l�O��|9�g3Q����s�`����R�tZ{�S�����~�'@����NC�'�4y<{���5�����?�n�>t���p����Q֕�߿�����񙦙˗� ��޽;F+`�����S*�4�%��9��Fw�Ǉ,��3K��glݽ;n�e��k�� ��dl������3d�qZ��Jѕ�H*�n*/}������؊�����mv�fܹ�g�{*,��qA�C���#�SM�v�|�&N;9)���O�!������l�w�m������O�P=Q`���a�w�����vo�����y�����S�o�˙��%��������l��:��"�X*ni���L�����k#l<\�n�G��Ҷ���E_�ȶKV�E��7�o��v��J;y�lYz+�S��:;x���+nD����A�ݏe"�]A�y���uWH֓N���{T U:Ur&W�nv2|���oє'��б#���u�7�����0h^T �x��ׯW���,׹�ᬭc�ScD��M��i4��`�C�`-����.r��:;ew������VN�I���h*_ďb�@e�����s�ι(0���(�X�J8$��YۅǏ��J�<��=y�dw����Wm�M���.��E�������!:Plp0W?��#�a^�����`W�}�p����4�\�Nɤ@
���=r��/�eU��a�?������������\���a��<���ə�K:�NC:�AAث}���AEᤤ��å�&	��%0��3�CT����z^2׌�܊�+�������{⭘L'�)Ҕ����|{� o3�0�Y���vX���+�=(�/CӨ��'����wT ����ö6��6� �,c:1(�C��,ȴ��;��9T�u �<ϳ�[Kdv�A�������)�A`IS^~c��涱| <�F�F��X{��o�B���xr�RtD��hݕU6mz �H��@�������?asK��UP���qj�a^؆���${ΣG�m,{�4�����g��g����7��PC��7��.igIl�[����^���)	]#���Z���ؔ�/��g��i��M�/�C��"�cSS%x�̑L3���x��Ѩ[OwBd����Y��v��H�HݚK�>�̞��/��;�؂��^�y���B&�E�!���2��	�-饸ɞx,�ɿ�X{�^{K�����G^ұ�I���d�����f�s�F���r����]�O�]:�*R�\0���H�[:z>��I��j#�Q�o�("zӡ�4 ��]�+1���{j�kW9�!h2�t\V�&��
t�.�x���M�ի����}d��0��*����Ύ���&&������(�i%:�7��v�d9��?�s�����)��ZHׅ�0)��b[��튅L�&��t��ԑ�wr}s%��M�""��dT��_T{������a��6����T.,$���E0/K6{��|�1�k��Μ���^�%3VPzb78n[g�:Uhn� �b�!�=�w=ō󤥽~���r������G��\��O�1mż������6�N���A����N�/S�o+n<�>@�}�B�yv'��"O�g���yV����<w�[}Ƕ=�X����6�[��s^�跔iu���osw�����c+Ģj��\��7y��e��e����Y�{� 0?�����ؗ���j	��v�[���Z�é��ffQ�B��r�I��]��LU3�,O�[��H�o�t�Ǳ�-Bṣ���l�����8A�ePW���,� yC���g�5�(o�>��x�V��rְ��`�k#��7:~��h�ǲ^���~-�(��-�� X��,�-}ȝl����3~�L�����G�}��oTk ���x�����˸A��g����r�E��=���֮� ����B�~/�Y-���mhh�Myzyy�~jl�d���H)���������ϭ�����~Z �r�옳&E�γ��W�՟�n��%B���FW���$����v@�>%�eo����`#�o�1{������}?ڄ÷(EW�
1���د�bժU�AY�S�3�d�=�h�`�?g�s�m��T�}����[����Q�@��X�M8d�?���l�P���VB3]&<�`�F�����m_�/>-�tG ܏?�[+�Q����]ʙ��4�Y�<���YAr5^�!��ΕV�oZ����|9p����a����ޯ�q�/�-�c��\����^�%��p��ٰ���yv�}E���rk�E�&e��v!�x��h)6������FTE+���R��T~̎2��c�{v�Cߝ���=��^���c_r��q��_8�P�}c�m����tkJ�I�A 殗W@m�2�Q�>=�y���������S�Qu=�P$�wO��^�R�V6"Nڗ�BŨk�V<9�r��}�~V�5�R/�g1���x����Ӛ�}daٶي�'��\������t4�k^˲&S ї~�2���+z���2UUU�6>�9�2)r�E�K&V	$�rǫߊC��hs���J�f�҅�=�6�P&tI�;�����1�����;��ڏ��F�1�����Cc4Y�O�ת���!,,��֡<����1���q\�)ļ"\GG:���!%���|���wo�����Mx�b��"?Ȕ��j��a+/\� p�b��oF[��FM��9y	�݉��b7-����בq_ԟg@�tS�pӺn�s�E�2[`Ai��V�R����.t�~��q�q�K`'�����J�e����kl�M,'���~Y�e���2��T��L�p���~]WwÕ݂��|٧})
J��ܗl��n����s��y����I&J�G3N�o�XOٻ#�Q��C`X���D	���ܬaВ�+PI^��7�]H�2<�}�X���k�7��c�1��	g!h�kF4GO�8v l4�2!�ѧ�Aڂ|��ؘ~�W~~�n)B�bD�$�Î�0߼V��v�b%"g������qGe��!f���|�$uP�&i��z�ze�Cs0X������T��<B��jM>{?^�a�Ĳ&<񈓟����0�#��]�n��W�'O����2���1�v�Z��J���V���4�z��"7'GGC%i4Ҁ]�wn���#���pȮ��������Yq��l��S��L�O~��[�BUx��D�wIl���`��K�D���s�Sw
3���W��W���?�?�w4���ʶ3>��K���^�0�M�j���=f�8j�A�D$�9��� &v��J��N��\�n��T���h�<<<�}w���A�_�h56�+.�G.�p-�6Q2:*@<x�X��A�+A�����^\/
䥉�X>���Շ��g=J�� ����k��bw
��ys`@��WD3�"�?y�d88g�Xs���̌�W�@6��qݕ�� %�.(�kxz��o�׭��۫QW��]5�zј'�H�c{�E�j�	A�l.��> -i�o�(Kq���d��XA�.����RZ�2͕o���0)��1��p��o��c�4qzd:)5u�z�)��G�UE֣0�O�������S�?~(��n_^�QE��Zy�Um�5xmii�F0%Ү)ۺJأ+��r!;V↸���R%�;��߯�����%m�Jz/�@Z8}yJ�������l�^?V��qo���_d���O++�ǁ��.bhE\7�rc�@u�敧?��Cml������$z��_%�d�0٥��|	}��~��U�1�,�	K�N��V��#W �B^�KN�I�B}��#��a\7�_2�M�sl!K�l��KG����bO��i6���K�rj|���-�cJ\�Oe}҆�e�����E��yk��--���n���WT�f漑���`p(y�IR9��C���G���`@�v7��"��؋3h�2 �C��
��Rf�B2کP�űw���_P�Ikn�y�����F	�Ϟ=��!��5 DP�jj*�9)ƫ����r�%��F�+,4��/ hv�>c�S�0��K���2c�����p��lc�%3�����9���3L#�-��]m<�%��ؾ4	"P�����4qڳ�wl2��ί��*��~r2�3�� �r_Ӣ���j�nYD�2� &��VMM�?�@��R�3��T��L�8��/6ō]�xi��rUܿ�:�1a!U�m�=��JP.����m"����8�ƍ��g����,r\��q'��lEo}�Js)��K�ĂR���s$~�CZ��+W�Va� v��aB4��{��om͈=p�=�[v�S�������"��c>�9�ջt�֛�W����
>>>@�A�T��bj���4�¯�M��0,*J�����i=�q�y��/���+?��W �62���-> >c�Ǳ��0u��b�KݹB[��)�t%#�z�.N%���m����$Ba<�1��1	u�O�܅M�T��'�rt�I^%a��MV </o#A�-4�:^Vyh��e��(� rLLLt��Kl\AI0�Z���B�7�?����#�g�'����!R�4�*� �EDD {�ת8U�	�j<�u�����AV��k֟m���+@tsg���ۧ�ѣG�I�T@���Y_��+�!P�S�}�ٛ����͉$Ā�U�����L"�hWm����T�:�^GQ�gN����V��:�����قDo分6ħ������P�e �W�W��i�=)���"*�aY}��<Lb��+Íe��.M��՜��_�p�sު�#�\�J���3	��b���dy�-��� �м��x�O=���-��_�)M��N�A��'h^C��B�qCLw��P.vlX��XL)U$��3���fbS�C�M�N͚y���1���#�����})������&�Nd:���-UtA��	�s�ǔf�f�X�3샠��ǔޟ�x�|���e��i�p�^�)Ps�+�[F>K.أ����$��'�璍��I�X�(M3��!Z��5}>Nb!�#�L7/7�/�|\l_��E�E� �2KZ�*����)�%�Ut�V�JDd�O�evv�����'��ڣk`Mސ̖����O�Q"��虦T�zM'f�����;!��4[*f懀��p�9 � �+w�c���o���%��Yh-Q�}�=�wCd��s��D��wlt�FRj��h��#)���;e*�J""�8�����F��O��~��x�` ޚ^�Fx�@��X_&�[k��_[KѶ��8������N��!i��ǎm��Q�X;��S]O�lP�!(k�f�*6���������w����v�����:������hc���B�=e��b����|���	\JJx_����!��/b��R!"�ѷ���hc�J=Q�!���9{�p�֭p -�?"w���齏d�n��\��8��\	�_nF��kqk�$�>���� 1q�b��jl�x�
�Nъ��k�������~�}�	`��
���伢�h�z��b&�t��"�++ɐ���!�E�d{.�;Ē�����8����B����M|�޽�������L�k�*߶x��Ծ"@^���kY+k�r8n��q0U�kl�#D��kF�m@��<R8�x��m�H�J������q;��R�9��ʝp���X&�Gؖ^��z�R����?p�ۣ���s�ӓ2U?�A���L���| b
ne,ie�㸪&���HV��;S�h��(�J����l��e����:wG�uq�D9CW��1�l��'��j�����~�o���$A=����5R��TV�Z!Bj8f��=��K��|=k�03���O���Q�I�V"�^��m��7�7�!�u�[��'UbN� ��8�=���i�~AFZ,��������~s/�OҐx>�9�'�dr����d�p��B��ߕSS%8������
��摚��C �u�-QKs�oo���t���CJf%)��W$�èΝ{v.��Dg+�8����cW�Ud,A�j<�	n�fU[�تN�j�ۨ�V�/M/���_A�8�Ly垊3y��\���ר
[�����ac�9��!9kH��f�
��a,����O�>��Q�/� ������ߴ��@!�� �Ii��nє�~4��S
D϶���1���r����d4̿Y,����h}��}X.�ζ��P�t�_��O]��3ܛ���a��ϚcJ�U�+�����k���X�&��m� �f��f�����g��N���g�M��[��n��	�,��#�"��²}�q���y!����#��~�u�ZRс�:X>[���+���o�.3P��m���N��1�P l��;7طXS�2�ס���/L�a�wV����$q20���W�F�@������loIE���Y��`}D��cx���\��T�W>�kPN�rS�����Yq��:�&���;O�cK��>�.ƚ[��+�;!*�mᔾ���ѕ[o���"d���P xHf=��z.@�Yb9ϸ�&�_�����Q��A@�S�А�|xBRo�F�EΙui(a:&F�րV�;{q*�������jx"��s5�e���'��[]��q��	�o��X�F]=-�)������R����	0�D��FY�!WG���'�Am��ϖ^;��c����OގmT��N\E��]*vU�7_�RM�T��3�:�Ҙ�M<�f&S;D;���Or ��j�1�M�P����
Dq��޺�5A�������A��$��دH
'���u���|�J^�u�iJY8�)<S�"��"D��A������LR���ou�^6�2x*�p����|6���~=�9q�l�?�>�i��.r��i�r��^�؈ٺ�H�1A8Hf�M(����I�V��u�Uw���]������O:(O�]$C�E �����wB/�3�{��m�#ߞ�<u��1�=�O��
$ݒ�C����Rԁ�`Wy�����M���h9} (�[��I����b7�a�l�t�+͟�� I� w�JJ�O���m��
'`)t
W����jQ��_�@ﮎe��u$����V�e�&mm5��f&���_ M�ț�IY&D�0�)�7��&^��!͟8;I�~�6�y�̺*̖��E��-]��|��:.Y���\����O���zzb,�>�?e�O��3#[f���;�YEn�F�d�}��:G<�y��?� ������B���޽��Dׅ�dve�~%@���5h)������7�ߠ\��|�`�����
�-V �ylso8��}:�Z�|�i�k1!�H�}�b>��e8u[��˳33�W�yL�w@a�O�����!l�AݙG0�rf܀�e�f|��	���`|ۼ����K��<���Zh-`c�������H�L�#�+h2Fl����D�=r����N`Z	MM�:r����Z���ڞ��k#�5��D�U̭�f��-Wn=�Ē#��d��%�T"T�w{��5ɴ���ǵ6����XF�xY��貘����n��;p,T��e��3S���X;����v-�V�uu��.��q���ByvU��Eb���Q��0A��Ӯˀ
����_*L3:z�z���)���}s��Z�%g��[���]D��N1�0	��T�f'���,c{�d�tښ��Q=���,;�u������9��-2iz��]� r'Ϟ�¼I(�7��/_��wp��N�B)��z%��M��W��t���tR��ڋ�R���5��ڍ�JOd-7lZ|E;W��w�8���H�Pٸ���g,�c]x�j�s��KAl!��`�1WY�&����Ӄ~��p��Q,��Nځo� ߒ�-8�D��	����Jtd�rJk�Hc'�2�K*�~�pGY�:�!<J��>SKz�3AI���=�������'�\>�MrR�U����|�N��}�����&uu����KΎW����E���W�/V`������L�d�𒂫��?��~�:��޿(5�F��tv8\7)T��8�z�O�6E�@F���-i�V.�f
n����YUE�j\Ai�?�2�0��2��߽�5��D�5�E�@��4l��@V�$�o�>���냅&�>Z��,��n��~�����C��H�D#�O����;�4g$<A��g䌍����G,v�j��v�H�c�,���ʥ�b� �-��<�фNC�aL�FSSI�w�r��vM&�����b9���Ր08�<��:68��������ߪ$Lߎ��B6��b��ԩ�Λ�8��ܹG%���2|ݕ�������/wet:M�TZ� &�bj�66'?���g�m�mw�xxxJ��Zz����O
��g�k����J��:oZ�`/�Dp�Q��g��}尢h�+//���X[+W�H��}'��O�tc"��X3�e>��$Ď����_�h�9��Y?'�2��4��Y�D�P�)/	t}s� $j_��X���=�P������ҫx���z�N������!����$����kb���B�}enϏu�R6�I�ιJxgRu�>$߬�,yJZ���2F��}�U����֯7PK]!�m�;߮�jY�����M�[�������,-�>l\��bԕ"�DG�u+;A=��O�I���|����tl����D���^�O`1��-X��s��7{�+��b8��Qn�ɧ�Ÿ��)*+�N6.��8�nx7VO���\s�r����`:�iee�E+^���)�H�^<18>��y57������#`�5np�/�M$�� ��S�������GK��Ϋ'�Tf+~���w����R�Z�7�]����*��2_|�s_��7�����w�n�#�{�L�=+ 2H/q�wu�C���=oK{�8�����HAv���	Xb�=b��)�~^c�e$(��T�����O��n��W�8���i|r:I��G-�yc�\k�N�f;u�"q�
�KԽ�.���ϗ~(��zO`��`|z���g�.��Њ�*�@���|@v����C	��T3�Ԇ9�l�>�l�f#(�8� v�'�h>�y�j�;q�&�]ˉG �]v��CТ�N��xz��+�r����6������SXtB��M��}�eY��=�gRʥ��	�as�j^/�VM!U_W=Q	���r�s�=xmt_}&�:��q\���&xE|�R,�.��W��o��ٸ�bW-C��T��&&x��Rʗb�q�c������+(�i�m���
��![)��#ɸ��>�Qr��k	L�����= h��,���z�?�m��}���Ên�R��81ԝ*��2dv���ߜ��!7�j�mj$ȍvj�G���s|��)Ǒ��T�W�z��������!O��vqMoC2q�η�$�Y-�n��{vZ-*`��v���ܛ�Py[Ww�lB�M"�̑�.'�����t[h��,R%�ƎC�C�z�陱r������<�f/4�+F����4��3�T�*u�p�y�c���*�&�*,M�ә���8߉���LO��{|��л̫o�w.��P�Ԑ�,`�ZZV]�#qY��W)*�h)����B�Y��gp���|���b�,n��7�\L�9�8X�(�e�Qn������G�Va-7��61�s8��<F?�=�����-t�
�W�� v,-pE{Y,y'9u��̔Ǌ���ew<�a�;��\������E�x�� Y���"K�v 
���˅��r|&]��L���#���+Wv�� ��Hݟ�0?,�Rـc�E�枀o�̃�kS͸�:�^	�i���#���e>���l��&8J��
��K6�g�`T�"�.y�(ث1�^���Gtx��2�vQ�H9� 5��1mS��L4�@�	~q�nR�j��ؕ���Y<ee���J:$����ݗ_��	�߾����&���.���_w(ߚ���Zo^YvȦ6���@E����(lMz%�y���˧��T�/�e��%�Ӂc� ���ʲ����(�q���3Jئ\2�͇+���+晼�L����������a��C�)2PY�^��spgf�-��F��S2�r1�`�®�����on��A~Tv�3��^~cSw��̉�G��E���h��?o�Fjٔ���	���NZZnuhN�ej� 4I�K��3 _�d����åƱ4��v�ƨ1Ww齁��j;.L�yy<Lɻ�[P���rqAE�#�c<��x(0�,;	1,��Bb>!�u�&�@���q�п08�C�c��F]Y�h��L�E��"4/)-
�Ѣw�&(�/���W\ė@��Fas��8<�H�f��?wӨ+?��+���8LMM�%���i#� ����D9��~�v�|�x�y�3,nU��1R05�854���"��/A��Y���.L3��#�\q��;�>�y'�s'qTV ���X�|59|�BMW�\����{����xߣgb�#���6C`���� ��	��|M
�����`Q_#9ە��>�� n�vE�G����޿��_=I�o;mD���_��։B����R�N<����s���,v��u��9LjП"Z�1�G�Y[;;ｩ���	`ݒ �0�&J#�;�?牿N|R@L�ŭ]���hۘ#�Uh�"��0�ڞξ��B3)q?@n����r�Z�!��/���Am� k�/P�#����սcc��5��d��,��]1�P�ae�z�� �T���4L70̂ �w0P��-�%d������K~�S+K%
}��~4pa���;��A��@�z��pn�R"���qia�Z3?�
W�Q6#��)L�^CQ�B���7�p���ʷF���j�7?>)�*��7z�Ƭ�����YiO��/���$���#�O���ۚ�&9;vf�=HM]1��0aEÞ�8|��G!0�d���]������.,�_�8�'XI˩��j���6zt�|�����K�����PIFtX���
�>��I��F�����J��%
8��}�&t����yD�0A�NZ� ����I�g��cVO0�����#��Ӄ��ŶI����c�o�ߐ�7}�4�!���o+N)���?�^��h���弍�U��e�g_q����X���I�I�$ 6*�-u}9{|�,�C���U������}�r�LC�86ʝ�ZJ��#��{�D��i���YJ����������O>�FQ�'eI��Gڅ>���d�"��s�Hc��r��/��r��'7یM߶|i����5�i5�lD���hXԝB�l�5[@��A}�/�"��u�RT`~x�	P6�����[9��8��o�ۈ6����w�$\/����y�r���
oh��m�n���qN�#RWw+
��I���Om;acC�I� y����b�!��i���l���dS��1)������T�Gۀ�	�u}.�r��j�?��g�]=�BBbdj��Đ��%��,��JNV٘��lR8���}R��-�l;������#�D���c/�wZ���p��V�A@<C���g���Y���y�������7��*��[�cfQ������8i�U�hlYË����E:s}�y��\
{>��[~\��~����d������ʥ�X�H{��������w��i,��� a�y�x���L��#0`A��yt���\»Oy�2�bt� �f;0ezs�t���b�?���������_c�*-!�e�ɂQ�4�E�K���b�j#�u`�Y5񈝷����=U@��]NK��~4���[ww�)|��ܼ��`���Ů�_=�����8-u�Z���^�N�L&����@��+���`>�dהl)J.(Z���c��Ж
G�pn辰�voX�Z����f���|y"A���w��x�L/}��m,m�C� N�m�Pf��}9�J���~ŭ=ئ�ŃG���{���G����j��Ñ�d���w�y��F���
AXH*U~��ˬ��gr�s�{n�FFF~�M����7��������qxv�es#�)�0PgF�7έ��|/�?���|܌�;�QC0h�3a~<@244�V>�����{�	e7(����?����^��-;ޔ��;���{D!����h>as"��������B��ٵѾz2�+5<�Y�_�+�Qhc�SC�qw'~����xLb,S�vтg}x�Z�
X�%�-�H��%��w����F:!99�|L5�i(�Rmc˯`��U}���k_�������o���Fe�ο���#g�6�k�6�'��ޙzˑ�Q����/����)����V͞S�����#������|P%��?��ݤ^��-���6Gc��a��=�`�.۷oy��Z��2��Y���V�Ë	�B����(��t�ҥG���Έ�����	�5'��M��8v���U!�ãf�/ (��(f&��>��'��7`i����b�s=��A��>@"5�[5�"@�LmR��-`!��ugp׬m%�Rd�<�A}�ѺDY��jk�=?����<��%�������?{�2�ʶk���JAW�u`����T��3����[�3���\֟B���˻�Y6���CoTktJ����[��~��;�#�����z|���ս%a�� ,Ȧ��Sd3�(J9���Q<�V09P\x��ף�T
����-֜<��IQhrhͭ�jb��V��F�롒�-QkB�|ݩ�t�)��!hSA�v���d[6V�Ib�IJ0�AKǃ,�C����i����m���b`��!R��3�8��;8���PDT���M�6�qꐑ�7P���N<�}x���-x���e�*@���;,��	�T�3��j���VkV`�n
"�9>L�w;Y���xj-��Ё�'�ͷ�\gr�N���(Ur�6�<�1�^����\8�|�X��+������/�8gn�������\�Xӯ���E&0I������?�bDeӼ�E��?������Y�K�6�ɨ�����0�2H:�[n?,�w�����V�c��w:�a��erl���
gc"5����|	���#_��o��ئ&�G����S?SW`�[�^���ԞYGn�G�]���e�L�m�ܣ�^cgq�����
RW�.%�{��=3��{�� ��5��M3�$O��H=�b��ע������F��W/�dB���V�Ӷ\����hir���6d�1�-�����£mUUU?��� A��9�}��O�._�����w(so�^i����� ��j
bħ(���w0Ֆ�0�jdve�x}�lG7%�Jh�%2��X�T�<�S�qQ{五g*�u����(���� ?���I��=W�n5��}�%��a�p��1��pG���㩃e�jb�:t`��8t�Luu�g.��3z�ײM�`���R��GYM�o��*�t�H�=�lNѾ�uW6n���x�ȉ�:�<�$�aC:��)��Z��'���q�v`="mQˤ1���ߘ��w�X�@E�"q�H�TB�]%�`��d��a�2,��0XJ�ɍ�a�uU�����ܹS�L����3}� xA�8M"�����?����\~�dᦢ���a��>f�Fk��<�%×�� �1��WT�ۗe0�x�,P� 
���ɓ�`�O�}A~5�PKv��tj�@v'=r�n����P8=)�{�D�:�l��X$�Y�_y"t�(��-��e?���)^`?���U!!H��_|@��.9>��$�=|8mvة�	;���
a�����M��Ϧ��#d#J��
%�_����#ݎ#U�N������l_�b�����q5��qMgs�9|eƾ}�9��D�����|9�^�d�Ԋ�A��q�F���V�}��d��J�j��y)i�9!"�s˶|��Ϻ�s��9sBl��~�d�:ցW�����kvm�#y�� �yK Rx|�e��+��1�(�[��,8\iu�X�MX`�Rq�1�J�%%����o�d���F�����<��Q(�EP�7{�~E�z�k�=%p�e��r�q��M���i3��dbGD����5My��uHaʆ�2�{�ȑ��ɍ��7�]����O2�5\��6X(��t�5�M�
M��p���u�d�u�n�aÛ�=���d��E��@\	N�e� ����B�OѾ������R�\�"��h�p'�İ���۶t��0��W�(�=qH��� ,ꉅ��'+m<�:t�[���-{{b��U�Qiz<����rT5���!�Bx(�!j�� �L�`.�stG�Y�ݟ���0�\�O�RR6��	��^��ێ�%	p�J:x��	�Z�Vka%P�p-f�����5r�Y��q>H�_T�&<@�K=0U���԰�R3���}!�l�(/����d��b ��`���+� P�#V���;tdq%�/�:��f������5� 3Q� <e�Ηau�~zT���B��V2mt�����+m�~<^� 	Q� jΪ��zI.�mSF?�?ۼFS�:m(=��?�Mҷ��s3}�b�ӿ���B-f/^��}]n�8�F,p��I�9���������A��=��\�zZ�]{��c?�Z����<'�B`K��䢕�'}m���ZW�����`��f�~Vl����-E8Y�g��6hS��-�d��KE��RrEC��GՕ�S�}�QI�"���I���L)�'C$SJ��x"�+I�
Ir�I2sJRd(S22e�<�����ߧ繍����z�����ڒ�y���(c����gé�Hi�6>�<3���j����A�7��=R�Ch*����q�g���'��2�n�����ߏ��1_R�j;ي/ٹ{��C~��]!�ӵ���n�
�1�5֦�E3�j�3�5k`��|��N���[0I���?�<��R�&�a�ڢk�u����f�n�M6�ͬg����~~���uӫvK�7�6rƊf�<)�����m������K�����mX/��f���D!J�f���~?�x��;�C�t���X'��ql��(�}�͝�EIT\�}}�����SFf�_s�+�\�6����;�����6N���r95��°߿YV5e���Ho�S[Q�A9����E̔0�蘚څ9����o?ڛ=�XPΞ���q�Af�W�\�񁺯-V�K��arzaJ�b�cZd�6�|R�`�nOrT�2�������D?vR%���J�:�sL�O:���J_r쳿Fq��9��CQ��f=�7D� ��h��QĜ�����m���<�o<���,��h�C�f����}ƙ�~e	���'����,�)@Vذl� {��0�*ĕ����# ��K�2��m�ӏUl�$��ަ	�[MMm�k�dvd{ȯ�\
p�.�#®��QQa3dJ�l��mg5��m�(Q��Ѵ�+�X2<CA8`��	T4���@U����sb���c&�1w���K���;�dў�'�brq���
D�}�����p���������dX<�zq�sG�33�&�c"��o�������r �)�&t�K	�!�`ÃA�f�iQ��a�>c��H�߿&��]u�
�iƚ?󬢢�Dv0/E2��U�,^���FGU)��&R����NNp���o6���y���!��(�̞��h��F�e���d����@ִBqp�[ RaV�a�~��O���~�Xt8����Ƞ\B*۔?sl۸Tf+W�h��#���+�l_fN~
��U�})S#E��*��%�;�+��/���t �nQ�0u�qa���v�����4�Z�|��G`�Ga��55�~3�r�,zܕ1{_ͪ����l�/\�'�nɂf'�r�CT^�2 �� �%g�3��x��?۸�����R�x����i3�Zi{|�*̮��0#�YGFK���m��������^rD;���iV���`	N�ls�c�B&Zl�1�V5DM���:Q妇�U>,�x��<�����o��cv�T�39��X�"�9���x��1���b��٭:�`��!����]Չ�����o�{u�����������iQ[I�=]���c�uNը�������W[�����DJ���������l���(�R砠 �a�&��@�^	��s0>�?�D<!@�`I:�w
����lC�&E������5��q�wvәfi�Z�W�߉8���0� �$�x�^n�R���%����D/G��G���i�+�bVݾ|�<E��*�}�/�?q�ق�P4;�YIf� F5���pǌ��"��d��T0ޘ	��x���/��*c��������	�����7%t��Y�$O�U��$D_2Ė�a��ɠ����G������Bd����c%�zW\z�ց��ӷ�������Đ��*��<�}]JB���6o����M����}�Sx[
m�p��:�!`V���e�����W�̾�L���]��!�8[��&��7US�����bO_��,�Rr�l��74�<??�Lw���� ��:��,�u!�����!�r.��\�q�w��\�7���l�������u9DF���މ5��-�رcG�P�Т/5�Φ���N��L{�(J�vwN�b�81E��6q�%_:���m}�Zat��8�x����~�p��p��lxxOր:�k���٧_3���|:	1h8;C���k����e��u1�\;cUw{�|F-�Ga�@���N�^��Kt#�;�q���?��/��1��<�ni����b�a�Si1[' /�eh������/��y�������K�Z5�PR����i�	��Ig�n��}2oϤg�M���ڶ�o��{�t�&������ȁi9#$�l)����բy��'�̪rނQ�O�>����#�0�I@�[~�`�?�L>E������[$�[�Mo!�z��� lη�tb�E�?�i(�N����u� ����^��7���1��>�M,�0��1x@���,�E����kE�� o�%Hs���\/N�ie!�g��7���T��"��>�X\499U��$	+��s�^[��st�<֛�D��<��#P�7�f��/H��F�$Fu1�O�EqQÝ�Н��ޜ�l��v�F��d5���N��s��ou������K����3��5%i)`��4��i	�!2Ũ�vK��C��>��}���3�w��4�y(��� ƆN9\�'---�pK�L1s�aؔ��ga��iA�G��~d/��圛*X�6q��惖��
>�O����#��kFi�m�4��8���Zk��q*���:@E__�����]�ߘWDx���rX&�"4�jƟ�ҏ7��Y��eu���[���ﳤ--y�*|�dU�Ht�y>/�ʠ:P5�ּn���=D����x���Unt�P��(`��|@h���ys�?	ƙ�!9yEFx��ipR�C�KArݔ!��UZ�Q`��^^^qJ�&�����N���1DxR~Bf�ɐ,� �u[�$L���������Ei�#���z��jjNZ(>gm�&f��Ivd����lv�[g�][�%�����w{�\ڮI?ܔ��M@��8�S+-d6���-�6�R7�r�Cx��^m	84j�Jɵ��Dz������8�瞙�R2�0�k�?+W��Hd-c���Pt�<g)�L�*��������Q�rPQ[|�2%ؚ6���a
�s����� 2o���-6$n\\P�pкL��o �M)��o$ڃ�d"�X�|;6c���u��-�,}q(��d��9r�X�(Bś|�3$�>�6�/h�.a�.c���|��#RY�En܌F��>}:�\c0�����k�@���$3�^��8���47��,x��<�pz������Pq~_�� ������7�C����A��\���x)���UB1�e<xvg�p�(�{j^X������nf/���}���f+���������Y�WM�E�|j���C���g�S�'��_fe1��?0����]�;Ȗ���ad�@�m괕�/	2��&|� �|Q"��Z[�H����D�-��;�o��t��Aw�,[��֢<�d�M��k_�l�Elj�' ���c0�'v"����*�Ν�b?4\mb�e��hk�D��s�.��k�V���f^�ۑ�{q,t��FB���׮5���f��,��?~<����F0zc��-���D�#���"�Pk/�ڤ�[X��6	������|R�м�=�2�擵-<�����Fh��D �#���.��:O�S�4�Y��_ؠ�tYRP�����r	`�l<
k���"�ׯ_���[6��)�[�J�xY �Zs1-�Y�@�g�	�[mC6v7n|(ݳ�O=�\'(��D�����9�9�h$HueO���̓�945�7<z��>U"!��j��v��Y?m���F~��W��θ�S9���-�3�)m���`��]�"�tV�ԕ�������@ψWiAQQy�&s� �7��>��s�bfJ��E�}2i�%>�Y��0�~<�w�BBy��ޜ��j.�ܿ6�&��ciڀ^]���f�g�ŷ3N�Vƶ%<���aV94�d^�4���#$������;[�Gи�k���yg+A(��i>�	�qe�}ef�5�%A�?[�X!X`�$F��tu F�[�*xo�y���65\�Ǜ��+����ky_2�*��(��C�`d�۱*�G��\<��iQ�9-��5����/Q�-'
�@�s�E�,�0�s臲~ky�h�A�|4��\�܎f�I�躉��`�H�zT.A������VۓՕ�,��k䵳$\쟃��W.�cmϿ��JK8����l�w�>���0Ss�T,��8������O�%��+�OL��D�K��h��E�����ܳ��>��~����EkM6�/���c��@<��N�L$�K-7�{�^��&s4��W�����V��î��e*<�|!{�����ց� ���ǂm�QaH�	�2���~~$Eh*����<�����g���u�orjW�l2WX� �)P��փ�a���i���@�ޤ�y���:�n(XT�T�䄱.��}u����(��I�4��<ڍ2�qs�������2e.��I��
�pr����щ9l�,R�!$n��W�0�N\�ݠ?`OT��7}������!�!�'��Q��W.uL�ܺ�",�,�ȋK7p����k�=��$v��'�"Q��l���C��y�I����[0����?@X%�?,��P�1`T����Cq˸.�AP��},����9B}lz!0�=����s�qv��7�S6205Pu=��#񻔬fa��UvY#�}t͒���������A���'��Gm���h�c1h��ل���/,���桡��,1���g�u��6���H �Ӿ!X,���:��f��*�Vrr2�t�|k�������I��+�b�59ς��S��]�t����7f��������?�P����+����.�?'����ccW1G�p�s�sz��mDc�`_��u��bHO[	d���m�����<m(�X>H�}K��af���:q�?�����ߓ'������|��ph�'XMm�'�U��ɐm�`���v�.ť"Q��Y�=D�ߒ������/Yq�v��5&��Ԝi�\�yU�����C�wpryy.�˫����E?q��(M���FK߾��S"xH>_���释R�%�9=ͥ��%A��f���
Ϭ?z-Zq�h�l������0�v8U,λc/W߼���m�D���|~�x �n���J��ԍl.A�-��E��X�z�o.]j�Z��SdRk�"n��u�,����`�
D���)�M���A@R�#&9r�+y�I�kSk���,��;W�73i�����cE疊g�F4S.`��ҙ�a�T���+<���Փ�q�W0�Q�a��:���/w2�3`��+��so�+�<Z�(�T)��{����S��R86%���u{�^^�g���N��>��l��x�ܙ.x����G���%𯜑��#��\)ż|���{���E/��H��U�Z�d�`ڂ>�jj���)�����̔Dqz�X[x�2#���E{�?9�6�ŘiY�ŀl=����m�۰0��`�U��m�����q���"$���|l��\>Dg���LOD��#q�،�U	'���9�������&H�����p���"�4���-s$C��_���;���������H��C�L���&�V�#XK��܏ƒ��&6�螋�^�.~�������]j�8�����i���<3��7���^�������=�>E �4#gЉ��I�%�"E璙�X1��V+_^�2alXmCy�*e����������*����l�TC�r�1��1;�#����!��eא�T{v��/|�L���{}VeKZ�%Ix��)���b�]Z���"<@��xlㄛY=��~4ʖ`�2��t�dЭ۷�~�"�9��;��.W|����^��G�=��8��װk.���dLw&N�27���8���^��P���VT����Ó��;ql�����UD�V\���>�Be�'�x�a>G�
��:��f�,���Io&����#`����(in7a��iۮ��ق7��a��L��//�g�K�[3��6r4�;�� y�llll��/����j�9J�>�5� iJ2����W~���&���A~>c��J�Ɨ����+;��^�W�J��(����_�Mҙ��s5v�}%�����K���#\8teW�Y3E';4�ڛ&������9�^,h�w >��
�tn~���WV�x���1�0����y�#�öb�yXM�,D �����Q��w��G�g�@�H^��E�C�� ��6�J��j'���?��θ��� >[�z��1\5� ۖK甠r�׬�ɤ� �����S�>m��L�G!H�_��	�mF.b��(����:d$jL�H�F�m�N�|-T"j�-���l�`���&?�	��@XD�O/}�ӯ��3�d_�:��� ը��Kh,�M��֭�Ϙs��'�7�����]Tñƙ)c��/Ҹu�y�p�(��6_���\�&�#�����@��w�g�#՚�M�`��&=�,n����C�z��(����ˈA�}����+7*��v_�B��ѣx�N�e���[��Ɵ�;��?Q߫���OGl��j#���D�c���N��Z�AF��y�,���nu�hl���`�r5�v��U��O@9����b�
�Y�����G��^� 7#�����}}�nb���	J!j�5��l�@�E���&נi>G��O��N:�u����m�h�(,� -Jd�1-fZk�\EW�6���L�߂�>n���Z�yv�/�S���p�n&s�y�
A��0�ԕ����
�Ѳ���-��'gKz�΋w��?�i��7��go��� L��*U\�q���R�׉�Iipη$��������c#�p��tx2���ϝ�lWI���[JX�䣼�:O�Y�鶤K��0*�	.#����gn�~a)S���]T�Ic�[ɖ&,D�2X��ܙS��PX+�c�
�A&���ߙ&����ڽw�����É������3�u��4�pt4�/�elt�}/�C��y��Z��K3_�m��Q�}�jT陶�7&<�=�-���{��B8��_.�Q�BK�T���� ���˲��/Kݧ���Boр�4�|�P;�������;�}<�]Q���@̶�HN7��ȄAy�8h���29lD*Dl� s�<q��3S#Ck0��ˊ���ON.Q��J�|�/�*��28�c!�[)���R��v���(�����g�]65��ՍEy���:v>P(�����J����|���J�~�/���O>�/n�(�]TVF��0I1�%�EE�g&c����|1�iL�I�P�3,�Wb�vOu�^�J�E<t�c����nX�	\(���Yr�p��1����jֽ��C]�#��"+.�lmp�ԏJ^��4ˏ���Z6 ɯIg^�&�R N�� n�;.�׭k�M�V)�ܺ{k��V��?�e-u��1_��"t���rǪ� UX��%��f��"���ٿ�7�1 ,��\u�~�� ;�i�k�͈y?O貈&�#��"}��p������/d!�
E�-,�7�� $I��k�
V��@l�qk�:h���K�C�24�G��[D3��gRA��g�?�eK��Eܩ������w��h�`El��	OD��)d�����)���[nS.6LĂ��+�ȉ0�W�|���5�G�b!(�0g��x]|j������l��Ƒw���»�W-�g����Dʑ}!���a%��~>Y�}�i�y��s��7|M�Z������?���a}��%�4����&�e7n����-�D�awψ�G�/[Ы�ީ%��_:W:�Կb�X�kɋ��H�T�*�����$s���	p�¶��M}t�y^K�ð�95gH���@�d^��:���#:�5� 6.��5x�q��`��X���҄6G��mN�h���Ėk��(/��F�td[�h��\!;�r�ۏ�;�B����FF�ɱ
V.|�c!L����nNl�ђ�KNNn�A���Wj��~�VhpMHɗ�VF�n�?�.��)�,��{F���ٕ�d���sOz�P��2��]��%����ǰ)**�������NJ:p��O2} ߾?}LC�T4�z��ըr�..�O[����gڅr��g�����zA�|K�
����b'�z�F�*<{��cǎ���z96�@ ���׉�6���(��r<	��yy˰k�vHKG�����GݶrQ�����.�5�-��>u���q[��v�2�k����i����"���Z�(KOIDc�ʲe�`�N$�R߻x��H5�*��	���T�{���ITԁ8�D\f�������Nl��������px�縤ÿ��/�&I���������yT��~~��>�E���+7o�����bX,�_I�,���$W��~gQK�~}�+�7��ec�V���o�,�x{�D%^��l޹��:>N��<<v�l� ̢47��xB�u⊐��W�DaK4�:��F.���!�u�Z�W�_"�Qk�����1�!&�-�/����������J;�`K��?�+W��ةbᥛ���Xc�>>��N6�c+ׄ�׀�ð�������h��.g�$�r(##C�j#�Fҩ,�/ߚx��j뙅���m��{W?����4ﲆlgj��]L�}�w}�|>�������n	NFBI���������/����Ck����R�^Ϯ<���q+�������Ű�����[��P��ZP�^F�}�?�7&���HH��Rp,�٬��eS^�҃؇��fS���}{׮]���×�,k��7���Sd��}"1{�!�a!��i�I1x���;����|c��4����V����`��`���w��lZ���Q)\d������xzB\@�R&��->�B�:q��퓘���KO��>(�!��y�U8/p##3'x�G��<�y�у)~�1)))�����	N����M��Y_���u��M>ߤ^�pr�E)�8�����CP����Y����`4梦��H��[Y(�hSO||��)��QII۰��jW1K>i��\������g6N%0g����Ne%1�=�3�
���.�xY��9�!��Ǥ[�s�P��8z�r�ke�A����SW׏&�LGs ��#�	�L�ۋF��Jo�%�U=zwmjWj�T<	�*E�[AZ�{P�q9�>bɂG��SSS�lm珸��
#�Zn�G-d�X�׀��u�gV�"�42ҳ<��ϻ~��sPj��KG��6�"���lD\A0ےO��G�¿�~{]�it�����}&a��B�2T�4��}�6�H>j__*{�b�Wt�mwCv�H'��ă�x"���T{{���h��h�����Ûz�^�m�������k��7/�T�.� ��)��ˢ��m�����[��/}��F�[ζ�FB�o�-�`����a`����}��{�њ�~��@�g�'E��;�m;�z_{g�Ά{I0�{��}vȝ0D�$*�P��`��+im0�Z�[��X�uU:<��4����e2���0�m�I��y(���
q����t���9PO��ę�ᨐ ]"�wL��iP]�i&Z�딂�F`�����F~���;l��|���x��ŋj����;�����Ԋ��c��x �أ��	A��a�!�_�^49~n5��{��0�bT@DP���6�^^ܼ4D�`��~B�Y[F���+� ���N��x\<�%��b��v�����O����ΉƙҚ� ~�{�UVF�A�H�NK}���w$��"	~��۟ hw-�?��b]A%��ԻnnNh����$��<�(��{�뾬�L�S�D�*���|�1z�حO����+�VU�[���P�Ĕ@�}x�6�:�B��/o�M�=�YQ�ͷw�#�f���S�>޵c�Y�@G�����܄���K҆���:�0� U|ɂOcT��36i-�y��I��#Sߌ]�w?}�ѱE.	$
���^���Bzn��{�OOM��+��	b���mh\;���<����i{�?|��"ԕQ�IYG`�j-8h�����ÿjΐY�QI�#����^l�S �^�(�|4H�h��������tu��B,�c�X=h8M��j���~�B ���� .�I ��C��� �?Sk��S�>�"�w+��σc����wd3�ϧ�'�cV�^]��/�2��;�����ncSn]�����=��m�(��ν'ɂp��Ғ�E��-AY��}��:L��17��#�>�q	:�̎�Ɯe���9�����@j<|��ۛL߾C�k]��v7F*�xrD���]�+j]�9�֊g"a!c��
H�Y�E�;255X�p�{�i���tE�u��M���}?����|�qn\CC��z�!S�{���
l��Rj�9�b��)�&��:x&���X֖�_۳��N���۠�B�pڡ�EJ�`����Fln:��N��맨�
�)�H��m{S�����[��+=u�����/^���bI��l��Q��"�$aV���k�3{��& �o�T����,����/ f+**s����,����!a9'��m�2a��Ȇ{LR�4��BE֜a����0��~�q�`��������~�)�p�Q�:u*�f�ׯ1<��{Vݎ���ܧCY�{ fz�e+}��5��\ś�d��%�)� �K(�g:ͭ�SD�>��=�+�zK�%;9�(�- �a��JHH���cw�/7�q�ZM�I 
�J�  .5d��N�M����'w�)#&դ�b%���P圕n�Eb�܋C����Ǆ�_N8�p�
}���:0�b'��/��Ǐ��T��mLܬ̯���x����>�O��{�5�4�"v� ���j+���w/��S�:2�}B�n�j�pAh�K�t^	!��O�j^8vk	Ah��~�Sf�Nq`�@�Ν;��
��ׯ6lذCQ1X7����*������x)q��h��,�3�]�7����hlL���:�Y7�L(���z3�uj�������'�`XD\���w�n_�����΍��w�M��):x/Y��V�4#fQ��kC�-l��5L�6DĲoLc����}�:�12X�
o�4�%�2Nwk�YsPg�� ��X�kL��Kkn4�'��M�X�jC�z3��W�eP� �V�:�<���n��#�'�z$#!֬��f������:����p����9%%��<��UU'�?�lMB����r衶x~e�rX�����l�	��Y"9<��FB�X&����E�8`j-�c{�szsg�=녀�0$�x������BӅ��5��M�z��Oן|k���F�fEA��~�.숍:ԒD��	��^�2F�HX`ј�J�2ƶ�:1u���Dk�e��z�RE��n��i��C�sxGF�چ�����NN�_m���`Cr���ǳhD.JƟ�����Y�e�ã�&R1@
���g#��ڼ�V�Y����W;�>�o��s�g��ѳ�s�x}�l���`�*j�!����)�q�����������*�Uގ�
���/����t:#�����|K�!��j��/hCD0���G�0M�;)�cQ�����Ez���+�ccdl?~�>C	9M�Ͼ<�P�Fsz�����{s��>̡��Ͽ���lu�\��Y�ݾQ�u�uÙ���a�s�s���%#����w��  ^�=����]��^+�cl��|�]~2��~ҝ���Kǎ�p�Nl�$.!��5��)))��Օ<�2��]���]05u_�\+/?ד���Ռ���s�Aߚ�����'-��s�X��	GMOPmC����f1��ؼr�ťݳU��r�wk+�,{��qX�K�.=*�_P �V$Y���H�ȹ��o/A)m�E� �|\�� ���n�+�nI�W�"qz�=����,&�%?�,���ۚ�,Lr&�l�
��3�y��P�u���^��'�ggww��o�����rs-�`i���n�2��Oz?R��TC�>��������/�� f8~������-r�&6I��$�Ory���_�0�|���	
<���4��ݖ��۾���ӴfY�������O
�msq}�(��b.x����E���>q���,��H����ǒkًY�v���|]6:@4��,x���v<�f��c�raU�#��������o��'�{q�e�B����-��������ei`�f����6Ny��� K���e� č��t<�����a����g�!cRq�L%��O�.��M��,�a"tq�"GP�����l-7�Pl-��4�1 s�v����B�_������
�/�˺�{�̼�o��� ��q��Ra&���ea���L2�0⡬~Q��1��#�i�� �&,.\xP=�wxx��Z;Wy='''��{Uy���
M2	]⁪�H�C�
6�N�6�,<%�It�=�@m�%إ��^y���UJ�Ƕ3�2�Է��ί z7��N8�������V���'�v��ܟ�+��oᬈ���?�ߓH��'  PƤ����gHs�(=Ot�|���kr��\cp<)���`�0�|)�?�w���Q�M����A���$���������潾b�EL��V�e��f���i(�����Bwn
S'}��ނĞK��;ͲU+�+M���5Zv��L�{o#�F�o��f��<C���b��;w�g�Q��3��r�wf(�x�f/蘾,�wŻ_��ؠ��WfE������RJj����\UV�i8�����kԃ�^]KKK�X�5Kʀ�T~�|:�V�D��Lo���^O�d��-�����*'&�Qژs1�o圥+:�S��%�;+s�P�}0L�38�1%�W��AU���}PFJ��Y\;��Pڳ8�ue�Z��8&}Y(��R����,���7ω+�Df�����{�^��0:u+��ɱ��X��\
�M___U�L\z�I�&���]��]�����oo�=pe��8L"'���ML�ji(��ּ���=��J$j�677�o��P֯����f�Pޯ�Z_kkk[�Nt̮dka����~��&4�1!ơ�yN�P���SwJ5)�L�%ӿ��i�jU�5����95$�ѯ9�N� ��k����~�.SΗl�M2�j�Ъ��:9;[�`�wpH����t�8Z=�Ә�ye~�̂��l]U�Zkp��(]�j�Ku0���[;;�I�oA��~�Q��U����']�r���o����U:���ŷ�
wwυw�������ק���Y���Z+2v��ȱ�-R�N(Y�?�hh��tU)\�[6sU?"%`P���̰�N۵kW\nn���_�~ý���}^����o�D3��Ŝ��0r��ԙ&g���y��p|G�3g����Q��Xa����S�z@�ߴ�����2
�Fa[\q�G��y�d���06�q�����UY�XY�P���0�!)$�nCq���I�y���߇/ʦ�(v���N�'Ŗǎk�M��:99)H�O������$bO�%�L����̄����®��{��ɸ����Z��n��� )�P|7�tq�."ѭj%�U[�(5^3~n���	Ԯ@[/�i.��z��N(\���㚜l�Sz��"���E?�r��2���Xk0���.�=�Y^�~���D��w�r�g����e�ʁ�XV����Ek���õy�ׂ&B�'M���'��o.t�`H`�0��������d-f�hWOM��5[s*I�U�td��5K���؃�$��k@�����ΐ����\X%�1�0�+d�;��gW~l��\Rz�˳ya)7��(V�V�M��;�����䀯���;ė�񚺺��~Y�|����@���m���a�;�#�*�$���_�:{z^��7Ӻ_��
��#��a��KȃO��8,Ḥ���\N��;���W|�J
�����.MP~L��Z�{ �Bu�p[Ϛĵ��%*�(Xrў��C�0�I�[m]�YO Ǒ�� a�sd��g?������� ��%1��`�~����U�*�S���AGT0	j���?<thPPZ�Fa��3���jr��6cڻ����9�=MX!�����/))���ءC��@7O'ǝf�_z��#�!�$���(Sxvj|����P5a�D���kS��gQmѹ��X���5,C7�Y>��?�7߉�r֋���Y�����K	hkh��;h���Ȁ/%%#���,B�|���~�U�%�U{��iB�N%�f���W�b�����.4T�f���?�]�>f�仵��������D��:q'6���|�+���z���-@U����xO$��}���>n�#Ye!������}u���ZH;��z��U�@Z��6���y2��T���hF�H\bb�[��tu�f��[\<<]���n"�����he�%�$/J��I�#�����ttG5����Oà�=��r�fB���o�*����6$8�E��"�g�6�n�yB��"#R�����Grc'ֿ`&n�^|�~��A�3�U�F��w�(m�`����4o���<.##H�yɯ��}��g��j���@��+^��E?��v7��A<'oci
��jقy��5�O�/���v�ϯg�OH��P�v�_~ɗ%1+�sJp.��/8�]���/������ghdĲ�G�"��N��ބ�PD��iF�e�2̡�9�ݜ��x�o��;��M� ��9��qꕏ�89w�t; ��!v5�[^�{�v{�N!,#�,����ru�b9���L�IF)��|b����%�H�KA�U �K������f��:\��<	�� ���-
:�N���� ���M=��A5�Y"v�h���ŏX5����2;w�0�<y�b�s����^�E������vwKۨ5f�x�DU�0J��_CH��_B��Sr���#�C�O</�u�Mѯ�c����{����>ڱ{�9�+R��o��-�1;���Ѡ�;C'��a����H���ߧD':�0�|4�U55W#;)b�ͦd��Y���_��*�?�u�6n�����ܿ��%��t�$�C=9ޕ�����p3���~�����5��}������(wWȁU;v,zp B2�o>��t�4ȴ'K��|n6��-���� ���m������|J7檦���/�����c��F5|Q٧�[�v�o�e�D��i]�ׯ_[uV��Y?v��=��~�.Y�|l��X�G`��T)����Im�s*@O��j*�1�"���m0�Є�-O"������5T}��K_���|E�[�_�9��ٛ��}s�(�4$,LG.���/?����l#��Us[�?C��/j��h�IK�[}9m��C�+��$�wt���/�_F{��!��q�h�ݰ؜����������ͻ�&� l��%�j�q�T�����	������:�B8�TS����r���0�;	�O��/��E<����6(��c��Gֲ��<w�ʸ�5 ��]��?/C���x4����{�w��ਫNYU*�ԑ�U��r�������M�X"P�>3U�R��F0�~|0zO<��zm�H����輛+/s�-.Ğ�?y���$,,����83IvDx� �sU�!�����H������y�mx��'�����4��ٽ��yb�7�e�f&R,*�w�Ej��Xv����k����؝�'�=�~���/���|���4*�@ww7,v����|�m�`�̡����s�����i�ov�q�����`y���9����V�2�-�}X[^��7�P8�\�H�GKr8سg����s�vp��Wb}��{�d���l�þ"�|����-���j2�إ�bxHCu��� ��y:תU�0�p���ӧ�Fd�m�A�S�;�|�����ѣ�d������&7��ec��si�:y�a�q��̗}��A �ݓ�b�vӹp)-�L "�5}n��~ �4)&.1G�������+qOC	���^�ܛ��_dp��A���Az+1�t��ID�^�f=p��Ҵ���с�mH�7��ft��ɾ���Ys���}M{q
ϵ��ݪ�����|C�ӧ�M�u�B��f/�K{��p������U`�w����8���Z�:�E����\(��]4�q,�7t�"G�+%g+:!9�\.⧵�<E	���Ź��Ҷr�F�`�V ����pQJ�T��#��c2eĘ�`eUͬ$1?�a敎o������c�N�]g_\�2����<W���w��UT<���.���=��������(�$�;wn����0:'����R!��/�/D��tD�c����+�ߢ,ү�8:��˱��rW��A���K"�D��\�s@�('�0�U����5�����	�|��(d�L��/M��,�蔛�`�H%�k�aI[���ʋk��66�k�Ld���Yt�IO?p_��з�q_GAXW.���'�R�M�s��!*'%&���#�s<����4\;��v�9�`��݇"(��J�؉X#�Ի[|fv�ܩ��%�m�T�5o��@����zW��χD*=��N��3n7�v����$f���2(��Q�}�E-�j2�@�y9�t�e�Z���(��jd�4LҫH͝�_�%��Q >���J'`w V��L�şJU�l�������R�<zIݬ�����p��΋_)U��ѨGg�H��W�(�87�8C� �&��'�cN��G�hU����T��x��(�+�K?}jטԈ�#��uMMk ����OOO/��*�T�_�2V);,@rn�xL���{�6%��m��<Q�~a���k9�w`�x-ʆ8��*��ϰ�j9��n�r��Z����@�3��'��K�p�18@}Xټ��Z �'����SY%͞n���?��֠S ��{MZ���|dbOf#�)S�M\u�{�����������p�L4Ú�չgf`OkF��d�L.
�'�0�0�/_�> �ohg�\��Mp��#a��c�,�wb�$&	�6X��l㞱#`����
�K7~C�V��3v 3qQЗ��������bը���ф�%{{m0�7&er��|��[���#s��r_���X*�k�=���sz@ԕ?z�v�uFD�Fu⡌e����xTѝژ��U���m|�A������[ �#�b"C��T�?~Ch([\��4/nU�n}��wː���2��~����ľ�G�
�'����KOOO���[==�aB�a3�N]��r%��]���z�G����.��%m��p��cAP��K����En�S��V�l��rX�P��C��Y,�#(���8i�x�),8a������s��5����n�q���*U���5\�݋��+@:}�Z���:/�4z��R�+�JJԑ\�z8')�q(����f{�3�.�h�����L#%��#*�|�q���L�UD�4̸��Eh��/*7�I�~� ���w&�������3��>=ћ��ƦR���|�W��E^�,.]J)�9���h�|�)Ї'�>��FV���_Q[��<��bej��Ӓ`,c�3�V��Ef�EVn�Դ�������속�m#G��0j�|~B�0|�L�A$D���Mi©��h�A`���.(ZpXo#A�B��o�9���o�|�XXH֚滒Ɖ5MR�R�? �����{`�|��=�p*,���i�������s�P����Ş�9��LKn��zk�N}����K[h�
�����	h�|x�}��xi�A�\c˪�I��Z�PMT����z��጗|���HhMo{��4�B+��k�Z���C*�/^Z�L�<�����b+7-<�����,��\/�-�NJ�RU�� b+�VD������M9謜^�4������!z����q��[�[F&H@��'P�-�r��ѭc�fWC��8�r+��4�� F��I����4ϛ�
%����zG�� �z;�ڏ{u!ؼ{�/|ͯ[�%eg���s)����Ӝ��c�8�~���؜\KR�o��9`zԬ���մ�Tڳ��7r	��Ũ��@�<ײ~<��솆�Ue6���Ƅ��r���kL���h��9Og�������:�/��.<Ml��wD[6���p���&w"3�߰�پ'�M<D�sr�td����7���4��V�
6�_������|L�>�u4���ï���:��R�-���\��c3��l%G��E~�1QQ^ZYUnN�:p�$Y�N������G��~��3 �����6���e`�y2�Ж�z{5���K <�N��Rߴ	��V�= ��<v��Yf�i~'��'5u�ίIg�V�Ц&F�N]�_����[�5��+H��B�����lj����w���g���@��~�:X�����]�2Ut��5�����d�Ӵ���X?�6�z����:�$pM��<4W�%��Z����s�� x�$=m&���.�7$��;~{i���
����L���|��k �J�>�	��/@�+�t����d�
����_��`��,H�i%y_Ē�+�%�ؤd��
���@�l�1��7%�8%
��K��ý�}<|Qq��x:
OH,��of�X6ʵ����A����5����b{-kE ����s+�iI&�Ĝ���T]ǋV	 ��~lt���W���n�-��u�%��IƳd%�I<�}����L�\ڽ������	�m��Ĥ	h���Mt(V�t/����Hw�*kg���c�\Cw͒�ώ���75��g,)�L�A�<"���H��v��si �]�v���
lE��-ك�� �cm�V�s�b�0�����۷X�y��wj|H�Յ */������`��(��J3tr�{}:��[����[ R���)��2�D+�l���w�-c;P�;��Km需�ӣ��t��I�?��j��,�/2����e�t��-���ҎEƣה��i<KM�E�C(����+�1��X�!���ޠs\�Gq#0�\
������2n�-��:����tk������81i�-��!t�2;Ya������6�=�m?Z� ����}AB�J (�g��N�����j�p��W
�X��X���ۻ>XF��rqP��W�����?݆�n�wpn�YsX���A�]&�!ec�q��⠋��]�уgc�@f:���S�?*�����
�?�rƑ����_��X��`��f�3~>#9���5�g�[�8�/~B��E��z�Rg��մX�t���d����~G�{}�_���y������@���_�iX��>�����:���mX��&���׺01-��<���SY�$uYGŖ9���c�:0P!�C�W�E��������H��;,�X�1x.,��(+�'%m�Z��B!��bA�_�xQ(��0�3�222Qظ��0~Ѣ��1���+��}dv��7vd_��e����>^�RmǤ10/�� �&��c0�G>E������g�>�/�:�Y����SzaD�@����m��}�N���ov5�]���팓�âf펵)��ygu@]77s����1���r6�_����wk}h�
����l?a(@�$��nKzo� �x`���@�����|�y�{є��"`��w]nٱ P�=��lqS��㉸<���;���o�
^_�yl�V#�����MZ1�����bE�y`Ǯ]������ⓒM���.�!bUϜY{�M��������/��ԃ^�	�lo��f�`;ʜ>�������¦������x}�?I�*0�H�P>��S����)��L�Y�p�|ŎپEx~�Eo���R��{1��V͖ó�t�[�e�����N���32� r�(]I�b-�����	\/L���xO��c�;�����~ь�'��[	��tX���t3��AE����}\�V���|��=�+�P9��B�;�{��P
O_ք����*��~�Kp�K5r
��Aue��)s�)�	�9���&VC�7���F:eP����c��l����.IQFIV�(��B�g����"��$��̒�23v���Y%	�{���|�������珞�}��u������\S�A�@"� n�.�fm`e���@�����ݩ�F�z�ÁU��y6���v>Kg��Np�-�2L�9Sd�(�ۏ�nl@�&�˼fZ�����@�d��阦a�ą8rOq�okOO�{Bc� �^�/��E�*�+ِH4���$B���C~��7i\/zL'��<������-@:��Oa�ԀqFjŮ0�A�ДNHc���=���ʼ�^����MSs>�XY5Dct������4Ľd��2}�1:#��h����VUUm8X39;ve���������h�2�g�Z󛳾d�4�"�l�K��8���͏x����p�4���y%�!����W|���{&�8�qą��li���$�����]�N���:�	�k���dE�4M�Mg�9�H1��kkm�:�m����U��q�@�t놦�Z���7x��4J�$�*��w��۽e���O��n�|����MWo��Sֶ�-��Y�HnJ�Z4?<aX�x눷�~4XY55k��yZÙ��r�L���&�w��M(�M'O��z R���L3l�iQ�QU��%�G�j�k�ب��/t+�S�����w�A"W���l�@=������Qj�I��H߿z������'�3�����}�1R��)�,*��!5F�ܟ8ti>!˪�;XE4���sa�T���?q�Z�F	붕��1p�
�j5�;"?����0Ae�:BO�v}q��?�����v���b�:㘄�����ŝu�żu*���*����M���'M�p1�>)�H�����w'$$�Q��xG�z��⤪�`�Q@p�S���r�ϜoJ�'�����N���[+����ӿ}��|��)�����̩�!�(7W��O��Ǯ.����İ�$�YE���FG/</,�m�����e�a��D��`�׭�\L���%�0�4"apz�)��g����(/O˶=�5l�)L90���Z�*�Ō��99j[��.K���<��!_��	D:���=�++F�|�%�ۀCg߿��E �"��n�eFr�������#�+�汑���D:@5k�.&K�(U�^?���%O����xE}J��ri�1S�ڰ��N���Ks�)/eoEE�\:"�9��0�"�x�	�Mx�%33S4�r?,����o���XU��2	���C�c� 팜���n�X%U�n����C�+1j��D*۸�E��!�N�7sxt>��c�b�{��VnzنU��s��U��s� Y��s����I�I��A�T�)
����Ѭ�j��@o�+�� ��N��~YG_?V�p��Le������g�^����i; -VxPurvz^�H�r7YV�� �Ѷ����$lى��|��.����g��=��h||<y�R�G����<������V/�����}����G�Đ�C*�)�o�N��YO�t�!OGW7���L� ��u��YO�&Էoۦ�ڻՆHU��TWAqR�kr{�>=U�;


`L|L`�KsCY�z�>�Fx�Mu�.%����lQ����"��N���I/��H��_�Q�3n�|sà����W�5!_
�cЗ��,u���-F�#���G'MF|�n���Q��J�{۾W�����=��3)���(���^-����)�W\����;���Ͳə�]�a�(K�rw"�@L�F�o� �Z)��'&�0��X���K/f��6'�w����U�*��C�����b$$S��e1)obb����![[<��ۻXw����
��w�q���L�@[���**d	�λ�������4���-�"nEO.Jo<�������Ғ�&�b��C���7���ۀ{j�y� K�.��ݴ�&w��{�Z9= ~2�geh�����e�A�$)<��ùE@ļ�ťщ����$��u��s��*��Ή�,L��`ڦ���<��~���7���Tm�j���+4������Z;�_�����
�R"ޝWM�t{w�==/�}�]`h8��Gc;/�����VH��ڞBY��� �GH��)x"�Xx��6NΨ��p4�$jO79��p�mt���bI�Rxl�<�L����t󑅪�fo߯'��as=��þQu4`�u�D�Ǐ�_�y�0Ģ��%���/n��($�y�r�4�o%9�tt�J<� �ىݣ�C	-x���I��G7T�/�l_8��Uқֶ��W��� � �?(.~_�����#���@�+��p�)�����5�Ƌ4����J<��6�%�9m����՘�m��c����*vh�@�2�_��Ϗ�8�+q}�╗Ig���ޝ���&�] �#�A���"�M3����iv�2��Eu���Ỗ��ay�%�����R�+j�
w��b��?�E�5Ƀ3WV.�m�vf���4��ѹ��[���%�3�)�x\�uwGG�Э])س����=)$m��N���s��43��˳�hX^{PBMKE�g��P#��J8���oыCڭ֍^-��Tr�����TZl	h[q�*m�.��Z�b���*V����C��'���_�8p�`ƃ��I�oR��9�x��1�	��.����C�KVXM##��V3��T�Xnc�����!�e��{���|R���RZl��.gf
b3�% y��]�ՋȨ�W��y��&o�i|]=�����%���C���ܼU���M�ʷ.l70�^��5AAA����TD\��l.pJ������	7Z�s�����8��(Mu��ѝx�0Ӏh������L5����*O�Omj#�3��-��#M���In`pΪ�De+'g��ԓ,^����/ܫ�RN	��*�8r0�xC�h�����C��g�������:|=�� �����@~WWW��%�u�����4z5�#z5A��,t�>�i�m��0P��(�g���l�T�l�j��Y��Su�d��y.�q >J|�Ǟ<x�`fv�ᑞ0�&�v��,�T���S��ae���	n� Tn���aFh\*���X�aq0�2[[g����r�Ae�;�	~�ׯ_�̴I��S�w�����{x⶧��e�����V�g�|��z��]D�ʧ<zYWw�E����~�浺���?'g�|@�Ф{�5�1�Qxt�_<�b�E
�d�4�<+[3��(	K{O��Fv��/۰�:��l������z��m۬gF[/8:͞'�5?:&�/��ڂ����0��M���w�u�$`�l{�t�����J��jeV> >؍Ç�}�}�otlL}�ʽ��ݨ�>v8V��Zn��^#��+!��/7�ϵ\D��S`��8�o�!nwG�s��W�i��@�!�H�f?��rV�� �9���:���䘋�����|����X�gv@�ƍ�~�[Q��Ω���qO�Rm�x���������xb�{BJmx��`�J�>����뒥�1fZ2���V�m�8pф�*��xn8i���}z��)�m�z�h��B��ZN_j����Yv]8���j����>[[[c	'���=�9b��kg,�x������oP�u�V��|1��.�Y��x؛fَ��VKcf���p����[lF�4d �VF
" ���,nq�U۹��h^�p�T�,a�B��3��
�w%��aU���E����x=�BCCC����&����u�6p"���b �����锱]rw�д�ٳG��ݔ���n��8�	>��S<D�66��?��&wKQ��Ϙ>�5�°~���;7����9��Ϳ<j���,jv��ݱq�0Ľ���˭0��t�*�34�|��Z�_���9�r���q3���6�iH,�*%�R�]13c�F����.Z����^���z7ڀ�s�_Y�O�����,���+�������%je||������[�&��?PH�V��kD��0��>RA��⌧�뇦S��� �������#��E�xt_�s<��,���@�=�"�Xک�Q����xfFF�ۍ4�;���r��cl?�w ^S�胻�o�yV���������{|�e��i����7��k����<:�� ���/b���>���U�*k �(�������ܰ(���1�#���17Nm#�,<kZz��W�5�Ϭ��?�KW���@t�~���,����eVD���Om�K���~�q*vv����nn��ꙴ
�7�������S�ab@rħ�����h�ä �)� 
������Q>�a�9�
��m��lg+���$1P��U��7eVF��x�����������H�LRCj�~�lI+Jk�9<�V���h�6�E�}G�R�B�!x'v$4�L"ه�w���/�����5.�N��9x( ������K�$9(� ��"�H����9p���X�=6 SRقj���JJZK'[K'I����m�1(���S���64X���3W�(��?�2��O�y0.��?�IxN1~��eB z�b��|�!�s�+�ω�HӜ�Z:KA��q����t�6�T矵IO������=1*��.]]�l���~^�Ml��� ���ǧ�4U�l��4��y���^& $,��=�� �3�����@�[ǹ��EN�oCl+黱�m0R?��,~�V�R���?�������!.q'6YI�јw����>}��E��5���!s
}��?<;��m�Tr�<:�3���7������\�ZX���1\:`ދ�ӕT��>?����>E��v�~O�����_/oV�$�^���h*�wwsN�ZL_4[:Af�B� ⸔ͷ��"z��:r��J�,G]SU���ZL` ���/�J����+�z ��|r��Bc�rwb��)�\��Q�99j���
��..Z��
���������2�x�^R"�;nk�li%j}�1)�U����MA��-�ed��բ���MF�s�x�Í^Y��>;�dT�۩�g;�Xq{-�
�����(�����4�FMؐ����D��|��.>����O//���¬���Z���Ol\�z\���d5R��X��;�dӰ�&��R��9c�MKߛ܆��l�>��i��|A����T^Q�H��al�Na��_����'�:��ʟķ7c�^���@�����`}�
T�uԔ	�I[����_���ey�7�i�K�����[��s�.�j�*]3��x{o����h��o����R�e<p�W�6}�3;�������I���5W�� �fKG���h��9�j����ɓ+�y�}Ea����mmm�wl[Vdl�� "�)��;��@ˉ��9377ھ#U�gq��9�pM���m�P�3`IK�8�KN�`g�U����{�+�%x��J�〒u9{���cc�Akc�-Ǆ�|,�z��X`-�����1��A�YI�U�ä Ģ}�SB	,�c��%��0^��i2��:�l��߬X�aYVbݾ8��b=�[Rb	{�)ŭ�S4x����]��0��kN������f�qRc����1.K��K��e6�g� �;::�֪��1S���s�x��6��(v�����j?��x��#������c<�0�V�ʮx��Q�����nn����|�>Y�gT�O�>e��L��6qy.ql:q����3���^ㅪVq�5�����\Ʌ����H�����n=���j�jGb�L�0?�6�0��Wn7� ��rr��^u��٩����&�N�NȽn�)s�k�4p�oM��`��l	'�cǎAt8�\� �ӓ3W/Nvg#D�����ϟ¨<V���X�ٸ�^#%�t���-���׹E�_��K��]~���!�U�VJ��j�@>��*��C���ؘ�`�h��]���UO}�Z��c%��WPP�HHF5is���L��f<��1c���U�CsC��3�f���_a��A�T%��"�q�q����d|�"�\f@5�>����~�'�.Q�3�ڇҀD?=�c�g�{��N�JeOC"?& �vG7d@X��^=<p
 lM`��t'mR�P��e1��4����8�%��x��j��|��B>���#^Eģ��ͪ�K{���W�&��P*�> ��Axޥc�4�Û���m�i��W$\on�:gm�ί��?�]�̶]���N��缽4�����#SWfV!�������Z���x�@0Dԝ��K�bJZe2�,<Շ�0~T�N�@�}���f�]CS�HSU2X�2VnQ�Q��1�q��ѿ6Ԁf���VW�0��*#�����=L�18����\��3�-�Ga���m��J�C7K/��HS���#�cF=�eT�*�Y��7�� $����J�/��8���� �[)�����y�6��u��|�C�c>��Hs�^�����k��7�E(�(�_�$R��}�'~L�����S��+G�o�<br�	ܬ�>r��ջ��w��c���w��P�m�)��L� �����u����soB&R���Y���=P����A?~L/(hs�~V74=:1�'-����Dl%�ͦ�=�t�DD6j�H]�w�:����f�wݤE����p�"h��~ɖ%)�(h�%r�i��J.�RdT.ҙ$o� �n���$�x�ד8��*<�� A��+[��Bڢ4?�gW����I��15*�k^I�J�A�#<$�4��0����X��P1VǗ��J&E��vG�?|xְ\8�fF�e�X�S�P�g��jg���	%u@��I��q��g;
P�[���Է���,���@��;Xr>1?O��>`�h7e�i�.a���w|_�V�����u,B��!p������M	�rF��i8أ��#�|�5w4?q�^�i6�v��6��Ei�����_��b�G�@��;!!Y�o���_����^�y��mFvI��V����]zV�qF�"�� xrsw��Pa�R�y�yH��@5�mzs�&D�{�wyƿ<?���d�o�i�����Go��}я�tF��[�[�TG&��^���Y����t�gzB>l��O�͙��6$6�6R���0�qw|��k� �����G�;!�Ԙ�����h��{bx�����4����T���l!�D0�j ��jZs`��R�an'���~�v*!����o@��(�-#!�i;ȳ��nL�i\��c��I}�����Ʃ�7n�"ֱ���.��-�2�^w.oX��	f^��]�NF��[���[6���V��#�^���m��T����<ˆ�%{�u�����^s�ɋ��=@�e�����!F�[5E�K�8EAT޲֊��wXI�H��Y�qUl����M�	q�<�#,0�&/~D6��DԜ�zO��m��M	J�ضm�!�Gs�mGN~H8���z�#Q'J�T2L�/���yr]�>Q�C��q`�=&�[���e#+������<"�T��"����*V�,i�T�o�N�6��Qa��zC�yUP�ęi*��VJa�iiiqR*0!�2�h.��A������{��P�d���v۝��ȟv�r�ؙܷ���67z�lɺ.o�:��v`k�w���؏���7���� ���	�th��`��z��A�߮��@���*�A��M;K3�8�γ�ȏXT���&�����գ���YD�U��~]���O^EG@�����z �.��6��_�p*.�2QU��D��t�C�(G�h��n�|ŵ�GE˩(��!�A����t0��7�`&��Hq�iń+o�o�e����eS���5�	�Miwr����C���~io'�E�� �I��8!��g�-ϥ��D����|~���W�Ew'U��{�� �>�Nb�L�P21�>� ���vǩ���tP�Q��0@ �u���p��O|e�?W7��UQI��d��r���t�x%�E1~�e�j<����t�X����Lov�"+��g�dbN�� ���|��� ���GĖR���q��<���;�����bW������+6-�h(�z8Ш�H�>3�nے�J#���_AQ�8w��YϮ7�dǌ4ĉ�_��ڭ���� 
����� �E�-k�#Txo;�R�> .~L{-Z�3�_1<X+#'m�?�ר h�7��1��p���G�SН;�+Y/� �/.Mc�)����x-(��d0�ӭ㩋��{:
�]�\��t�� ��?�jO���뱳r�3!�##/�#*�S��f+r�|4|]����^�L���3Xy��5�C5H�e�wȜ��Ws�aՁ��O�l.rZ'�H&890�~��/\���x�[���R dhd���cq����`�4���5]�e6�j<x`+�~�mf�jdi�HD���#~f+������8��V�����H���vw��T}K�d7�('K���0��L��E�ش��n-�*�@sP*��r:ٓ���R���˗�Z�:[P�Ha�l�����.E���(�������b:�iH5�����#��`��d"3��`h�ަ1N���`�t�Ǟ�B?�XQ0���5�֦�0��^!�69?@^���T�AK6Q_:^6ٿۙ`V^����C�6vvoݪ5��l����/����s�.�~=�u����P\�����DO�H�G�^�o�L	����O�!G�]D�Z��ȑ���g���e�|��X����6� �SȂ:;3�M�Æ�������G��	��|���vx�҈<���ߝ(_p��e�Lo&y��+r5��o���c��w{r����t6b�L�o�į����"�ސ�������y����dǹ������Q�_���s���5�-���R�{��w���b:�����5�A^�jd7����̭�������������U�8�ߑ�d��x�`�?q��$�?���4
�2���� �5���0������L��.��E�V%HJ%Y\�#�*z�FƉ����悤��W���<y[
X�j�B}�ƻ��� F��Pr���w��8��\L�1���<�o�$�dӊ��)��m��:�N���b&�	�uJc�?Ug�Y	{%� �wl�@�?�|׾�ŤpXM%#;����3B�
�g�QN��p�^/�hۉ�!8]�h�M�//l۾],�����0?<���jt�aXGMI�1�i'�;�tU����׻��h�x�\}�E��\K�E[_?���r�Ҙh��'�c �q�/A����T�w�� ��mF�#�b�ڲ�nOtSiL�.��Dg1ٹth�m�����|S/�;m/\ ����A�P�`�:N�D���3�R�
FjI�;+[��w�"^Gq*Zx�{��-;�FpF��G�K�T��j�6�$P^@y�U���h'ĉ@�߸�P�N�� P�H��.���~���ts|�����H26�	���3N?�����v�����]~�U�>����y5{�@b��YA��w/�P��׉�Ň����|�X��I4��ǜ��;wb% D����}~�jk��4l�u'�Z���p�Y����f�������5���b�s5Q���mLr}�r[�VZ)x�I���'��|ⷃ@�	F
��,��THFO��D���0{II�e���.�#������bw��_�Xb��i�_TZc' �+�q`��{�0(!k K(�Ec�;9I
���U�JD2J
X�)N_x��fp�[va��⡄�	��Z�C�r�v沲2X�8JX`gvE�i�^��9�Q��tK����Z�`��,����"����*i��99j79�0���"?��SD<NH��J@r���K�^E���R�\v�ش�W��lK�-�.�Ϩ(5������i��?��V��̮@�A~�X���,NG� ������3I��KIe(��g���?'�S�~}�͵��Mv<���)����� &���&!���܂~��[x�M�(P8ցmA�R��<�x�ϳ��?�~��@��F�9S����>A��\Z��/�����a�DC����F��1T��%DEQP��s�
�������;8C\�d0����O+g쾚�,
��������w�-�V���{��x�$N�=q���}�2�a)�On�9Y��x��BDuA�R22N���C͑�ɋ\�(K�<�R�}N<�������ĉ��e� �*��� \�z�r����;6�:��D�q���J�u׏ޗ��:����%B�B��$#55��A�����D�&D)XB�*�C|ȿ8p`�x��$�^	���u�G��3�����T�h:���[���t��E�������'�7�r����!�����sܪ�a�sl5/o�-�?a�u�H�1�`�\Q9�Ez����?t���Ļ��&�\�1�4<��:����5`=�##��b�x�y�^�ӧ�s>	�2"8R���5�u�hp?�~%W;t�J�"�����	�)M{b�	�� ӸҨ�0m����M�p��DŲ��]	OI���M������6�5+�;�~�Q%�\$����V
���ʷ�����A����x��~OI��G�
��70���%"�A�a��?�o��zS�9�u����!u^/OY��A{b�,�����oV�qe����Z��'��!����E�?��?�LO�pt��־��68�08=��F �ފ5�T��U'g��`���k�A�8��/�w����ֹ�D�W����?<���@��B�:��}2���^U���V��)�<�QS�t~�0�2�_@1^�����ת�@'U�p�?�1V������t%��pvͦ��}c��^�l<��Op\w�a��
�����5�8aDz�����y<ڄ��~i�qܔk�0�G�)��S�L�P=�U��|/u��!ȼbDC�of��]��TiiϟG�T��H6��Mt�X�_mc�w�\�M�k���6���uCӰ���m��%�d�
�4IZb (���^c�+��{��Gw�Z6Dŷ-�V~��֖��i3,�e�8�F�=��Ȥ��s~��4k�������_&"�!��2���/<��]}�"榖'��V��&J��_����Q�Ϩ@e(�{�my:��r�4�֬TL��ZD��>C>�fhZ �������~?�|HD&��s�$�=�a?v�*����QMKK��_$2�$1+"�<t�sp�ԸӶ�{,F��Jo�E�/��0�3/z��*,,L���XR+�-��'D�� ߠVzq���'ά�`������5n��6M	���"(p�w͎l+�]&	QKW[;|��"�2l��`һ9ؒX��j����B�pmm��~��C�(�v@��H������eK�c8rۉ�J�ɳI��8���IG)2-�b��#8A�☨�R`������M� jL�"���E�?�Z{��N��P��; ������u���������p��52!�tN4s88oe���AV%�R1�j]ks�~��P�)>̒��<]��G����<�`=$�����7˷T&�
>�5څH;p�QZ��rrr26������ׂ@��pl�Z���R�7�Php�dTR?�[����sv{q�/�ЧJ�|1�F��JojJ
FeJ{D�zC ��G���R�s?���H~m@Tٻ�h�&6{` �R�&������N�����Qf���'��2]=Ft�?p�Mm�E��_���:��wyxF542�����2���.��a� `�K�#X F8�p�)EK ��,����r��eX=Ķ���I� ��Z��:*a @&z5����vɨ�t�+��k\��7������/�J<g��&71����[�.f#��wp��%v�jR���.R���N�ˁ�1f��ŉ�^��l$�G��)��Ő8 wo[q�q�ڕ�+)�^Y~: 1���x���+�'&��]���V�����ssz�b�1iT�ԁv��Cj8��+%�w����)c���e=]��Um�7�a�b���"����A�}4�� ���;��w��)0#Z��*�5��Kn�⒀�GY
�*���!�2��e�/�����"�E��z_�1"��R<� !B�� _�d��Mc��Y6��s �_�j��������7�Sa���o�o�P�+��=��Jf���	�;{{�|���w�_?����*�M�1{��;0��G��v׮ى	�����/Q��qݿs�i3cjt
����d	����Y�%O�Ծ����m7�[�ur�O �O=�HL��s-�NƗ�姇����`��#�}ǌ���1&�9;v��ruU>Hoo�Zji`��B䗎����w��6+��i�/Jn�S{e^�5�T�␌��g�~j�!"n�Ig��8�Lx��7����epظ�����X���V�x��p�˫ ƽA���.��F؋�_�&��7��6��`!rrȎYXT͕�+鹁����p韏l=<
]��F�	�Uf�x��V����v����<������'����a��G"pi^������P����SgIp��
������J<��\�A�S����L�WU���m҈{�������B!�<22�|c�vX����/��AړD��~�b)��	�D�sPgHPGǗ/�����(
L/,3�8nr�a3�(�=�$01���5�̗�Ƚ	\�
"B��Bp-�(�7��&�S�Ͽ�o���]]]%,�$.��ڵ��\����#�"����D�!�+�2ʭ��Y5��=W��g�¼ɔPEO.b��2�$Cl$s�j|�[X98Z[�����M���	v�´2"8����ro7!�?!������a�Ma|#씰���¦�N��Ԡ	T�z%�aXj k a"�L֩�|��J�=<��dLK<�j{ O�����e�@�c��a!�o�|T�%ҡr������Ā8K�fe����R�����Gn�d� 1�L���9Q�vw������#��11޼tx;wm��t����k�M��~ a��Qes�b�+e[D���FT����Ux���w:�;�,�MR�]��ߊ=��]�A��h;ߵ�����1�*������ ��lْ��ʳ��RP-�h�^��� ���yl����Y��w��˘�#�>�Bʑ�
 �l��0�X=�w��c�wy0�hT[�O���4F:Z"�\�*��Alj����O��'[���)B��͛k�Tpj��w�.X[��HKK77�H��n�12^�#6q�:Ī	u��>[F��������N��aA\��n��u���%?+�B	>)���V����"!�9�k��rG�U�+;����:Yee��GH�&d�o�P���2 ��U�Ԡ���Ս`QMcz��7ٶ	a��Jb��hߍ�j��<	���<<��d}:3m��#+���ȕ��{bֹ���#"��������DD-�m���Ьc��#��IP��	�����5y?�X��#����76pH#�V�W�@C�����r� [<v9��~�� 37wHV"�
zte)�ް�su�r�_gZC�iɮqԸ]70��^��}��Vln}�E])�[Sb��~�p�/~����(��M5���ӛ666g#bBC7�w==�x�����8)ע���6�s���k��&�� ����C��Z�TV�?L�d�E��6@��`wpK�jfNN[g�kq�z|����K'G�X��ǹ<7y%y9&T�<��`�+T&ĕ]Uj$&�����<�;oSh8!�z���H�LAoY��ֵ���H�4�Uxwu0c=����[�n�+O�&}�oo5�CI�^����go�����5�g;~��ڵ�*_���^�u�������Xƛ�,��1<�|b���T���g�~��~�5gױ��n���1�gz�Q���g������2,[5�g;��o߾�@�G�ܦ��§~��h��b5<ZY�1�(+�&Z�䌌[�;V,=���b�Q�����OC���ϟ"̵��ji�3^�n����'bcc�W�L��}�e����[3��H�Ѻ�L`����s-k9"�8�ԟ<v��"'jtC���ۑq���r����C����%5�� 1P3Fw���N���U�!�`�;�|w���7����bc�ɲ�l���9�P�:OJ�t�����j���~E)�b����A�'�,��{�S4m�ι��8@4:��������$�1�;*�'	��G��皵��edp�oQ^؋:�8�q��"B�Wu�Hw�������G�3�b�+��4�l� ��Q{�!o�b)�	�4���ꝝ�[w�C�ld5��ǐ~'(h�ˣGW8��1^f�b��� �qr�����~ӱ=���� �OZ��& <��&w^;��Dlc%�q�M����g����>x�jU�����̭�?���FZ��^O
��-�������ASr�n�C�b�ؔ���ߣ����tny��ك��w��t���3�a�T �!#7�S�D�妡��������/ ?8M��r唁����D���SSO�9&6�\'+�C ��xI)'��ΐ�9Y�˱��zCCCP���P�+��W�x��Yz�Ntcg�y�o�*�ݸ��������*�h�\X4�-�+)�JB���2N|���*l"����W^n�9䀴�Pӑm�>~<^�e`M�ň�o�Γ�HEW!Rb_$����^e�&&d�%o7< Іك�y��_�&�SRv�K:�2k��|����b���䗊�ܒKөॺ���_�,��7x^P �l��/O-�f�4�k�9�mph���r&��v��$c�ղ�ס�$EG�P�L؊�јL���o� A�?Qkdl���e��ؖ��_�zK׺�z|컴KbL̙��<���>���\u��7��L�uc3�	oz >1��I�K[�[�W*�'����K8�'�޽}�^Qa�U�%%"�����Hf������ί���I.v��;"bq�Jb����22�FF��T�?<���ĕ�h�va���ܢ-���@D�nW!
\��5z-@Kh�/��+y]�^$7#Ә;�=��7�tb�)q(i3ё�{��V����f�������*�5T�wQ�c%	�<�b��;4��w5�����-`�:�#+�Έ�r;؅�C�{�w ��OO�>�:B��S����s\�\E._2ʹV>r�L�o|��D�q0�����m �=� �t�̀,�W	�`5�(V��@ �F��D���3E�?�.XD��=�Xlnn�����Cb��@g��x�l����o��T �رs������
ax�\u���%ba���p$66^�y�m�77�6���������q��MuKҕ����O���1�k�����y�E���`�g{ϟ�\r9(G����,������2ܼ��.��PN�b�`��=5
�4У؟O;��t�G�+"ē�7�EY��_s����a+9q�E�V��v���'����J̤�-���1ִ�J#�ׄߵ�ym��(А�_����^qR���Z��J<{z�����bP��F�q�<������d�0sD��ͳ�Q|��9�˵	�#��Q�Q�س^���f���{r�_�����p`�u���wV��W%�ͫH�>X愭^@j*/�@و��$X��T�*��ʐ��o���M"%o8 ��$;�D�ﶛ��99�e����cciy�b�k��gk'�'�=��I?#�V]�H�q�����x"C�=��z9!La��2��a���Ȧ���򅻤)^Re'"6� +�QQQ�z�Mq,��ߩc����Y3>�Z,�RSv�3إ�������Oהx^	,��U%&�B��� q�2�R`�p��j���@G�Q��%��n�mI]���O�>���f�8~�ؖ�\'%hua��CK1!֭`B��d�� ?O���#��$�ծ�	Og@��Iȳ���	��i�����*�al��y02b���M��u�_訞�F��|�^��o"���B��*uL�;m��S:^�x�Q��Ph4�VrV�D����ց�Gd���R<[�,||��*��@�aRYY��L����	�����}�Nk�42VLZ���D�&�!W�ݵ�cc��ce��]W[��f�6ĉ^r�ô�ps���gŌ)��heD��r��S�����4��9()ɟ۞51ွ:�0�ς�ܑ�~O��H9�V}G�k��/\���U�X�hc�c�{�E&qjiܡk��	AJ����>'�K�������#Ϥ�S��O�LqS:ׯ�`��[[~z���z�'�5�^F��_�d�,��>�}v��F|�egy0
���"_K�*7z'#�4m___�b�T�'kA��Z�#�?��،`��@��j�V�J�!�����^0r�6A|z48h/�k��V����{���
������~����49���"a���_��"�2<:��z���
X=v|P�XY��Y5������>[I��B����I���|���Ǚf�g�`�-�$D����G#H��ikB,b�z��W]�P�z<�	O������
�0�7�b>S��>`W�FFb�.M}q���*���>i�^4�u���
��J�/��bц �׍o���5x�1�����&����W��x����u�lG�\������;�A谓�a�̉Ā	K��Y�_A�t� �MC���eӍ2Hw��v��E�L7\�n��Xv�*�ףR&"G�nr����� �����o�蕃�m,���9F�l۠�C�2@���+ޡj���K��U�xB���|Y^�l�$:qf�i���Şe���lhh�b�������5��L�͖J{L�a]����/'G��!��������<b��ZZ���̈́�����x��ӣ���K��ю���|�{����A��֖���Y*���6�* ��1���7��7��>��g�j�-x�	���sXjlTS���*v��rh:�������L���)M;�_�8���J���.MBZ��
��s�k;�9wH�+�<3��]��ȕ[�kRNk�[�Z�ء'�B���rU�o+��ѳ�����Do�9Q6�e�58v���}r�=x����<kqr\qNKp�r=�o/�6���n���o���i�yEn(�0Բ��
DW��ѭ[k��i�L��Վ�}��#>9��;�}i�c��pfr�1�蘠Ը��ֆ7H�͏fa+�A��k�@^rb\h�����3e�;E�<�S���Ot����M�!��6"�`����Y͐�Z�.�%������FO$��}~,lV�����(�?����$�>y��w8�؜_/鸬�6v�ݤ˜�J���?�=�r{�K!V�����˪y$�k�?@�<�Ħ��V]$U�)za����+�����M	�HA&z<[�K�m���AT
�N��w{H�+������ӓ�K�$%��o���q)�紵��	&{�/ߡ�z���8w���G��2'3���j�����h�r8u'�#~~ة�Y��Df�WWnܸ�4K F%��7�=��Z�49ɍ�����@9kj�@0F傋KXx������?�~8����~���ZG���!:�ޠ�9�+ �%��}��y++<i�i	PJG����4�%�L.��O����	�w�<�a{��40 �"3�"9
�k���c�|���*�,�A���n�dS�Gmz�UߓC�!#D�#�<�J%:��s��rIvF0�=,�1\5R<9�� ��L�8ΐ7��� ��yzff�>���<ݴ8俔��8���I��&,-��U!�)P����f�ǽ�w����|�_������N:��I�[s�U�}�(��dç���a�c�[߭'*{p
����~1����e��p;�� ��*+�E�n�x?3�^̻�(|
Q�����ԋ/k9R��P?��adT��A2�/�� ���G)׎_�^#��;�@�J$��hLD�d4�JB��0�ߟ�~����X	�o��bۍ�RP?*�p�ҏ�}J_s��QWWWТy���d������ܐcZ�*��edR��o&W����[�0i��gd�gdR"�й�B�wWEOӭu��lٮ]��[��޺ϡ�5��#v	�M5�a�[�����߹i�!�D��7���޽�(-���o+������jGn�!�B�	�|����������?�3i��,�@�_�@n&z��w�tO��1���[5f���T��o֖-L����y{ˤ��T�#ј u�V�.�4�c���F3��oCCRu]`��� �W�� ��IR(��g I=i�@X�H�GJNl����<r�E%��(�ma7P�<�'M������΢��^�k�|�^�����oz;�<��g�Y�0�zP��E>��Zf����p�
q�,�x�|����r3ʀJ��~�b��R$yVUS\��7C�zdƄH
b��52ܜ��<�����j�T=D*��5rKO�=�כ���D�B�diܻwoF~~����Q`Պ-�`����07�x�7yB����a��\���ؿ������a����	4$*�e?~l^����˽�z=�g���,O���I�eo� Fs�"�&��,llNbzn!\���'��.H��Ȋ77Bs���P
?�+[ۃ+�\���)d��Q�'�&���������R<�yRKQ�.mc{��ܳ��
�G*���I����x3;�fe��*̚��^v������m�����v�.��Xi�����M��n�Ks =Ly��t��ɀD:1==�m۶8R �Εã����6��+r��f���eaa�Z_ۅ����zt[�ũ�T����u��@&�/���GvH��_��:��ô�&P���y��W�*�j( ������%��9��h�G��Q.u�e���>�w�{(��		��QY���\߸��w)�)NH8v�.u�����v���cy�r��+���t%��A������J<��N��P� ���q��m���C���x+zr�!��=�\nn�,�i3�kc$�������c^L[9uS��@�'��%�7���YI6���$���ݽ�Vfq�9y��}�-;s�U+����i�#Ԅ�:�F#���pʼ�?"q�h�%Vn{��
 ��X_�ZzGa��i�T��\ٜ���y`��@p?!��߿_yЃ( 3��g� \b�,⡳$�J+���ѕk�vl��hBT����X;�գ�� �.����Ļ�/֯$1�b���}�}�.�N`c��D�]Ξ=�f�����'��'�7}��L��]�&�|L3t�ݔ���V�
��� P���|���[� Nh�3����	���ib QO& ��o�|�@�&�兞vLr@��A��j1��]�{r�EV�
������r�WaX}#1��YYY�ͧ�* �F����̧&��0^�����>��;������_[��Uˠ��"�\KS7��?fٺku�~��6�4~�_�q���HK�y,GPG�Ug�p?}��f���.H`P���d�GGpwa�;��엓��X����� "Dⷶΰ$`S%�?v�L���f��sk�����k��+�`׬�Hzu�B� ?Щ��

�924��9Pp��.;� c�=ǣG(�<{��R�bS8
���pt�L�>5@/����S����@^�3�37���p^>�-�td�@ipgMM�a��t��SuZmKc.��-�?�8�F�L�\1�F��67� U�bc B�)J""�u���2og6\y���Ef�>�`���[��e��_F����2�$�Ւd��B"#{e�v�$;+y�$;�a'��M	%�m���u{���=޷�>���t_�u����|��̀�o���h,�;�Fř���2���L*����})�ݿ��)�29��ϟWs
��� �#�Ey��A��d���t$%�J����:�+Cͻ��D>!�����/�ı�8���(�$�J��64<���6�G菓O��B��ed_�)ǀ�� �#�^
�|-��2;#P����]��2B�c����b�3��_c0����T����.,��FƧk�3<���$�"$+����,.t-6}���(׽���.d,�"KJK/�[���c&��_ZB���ЦA]݈䔔��BK��K��636��s��C�ș��`��,F�?�_�f�:Gz�ӝUϜ9���4��첥�Cr� �����<���]~���F��c� �B˃��܄�M�l8��ޒ�~z<,2�-�pop~�k��&�����vlOiJ�fBZ����������kR��̜��R��!�G���0����Ғd�}F���C�_`c���罈f��C
�{��R����N��6�c+�Sn�(�T�]��q�}a!���=�*K��Y=�F�6b��ɀn���8F��>r�1����^���!�l��U��}R��ѕq���z�l* d�;��u���-�M��!��v	�zF;�)����o�V��q����h�R��ְl
�dW"��Cfffd4��^m��եK��~�x���(�󇲌�ꊪ�I�Kܝ�q�l �zLCmW�����͍����E��_��O�PR*y=?83����j���<0�p>9yy����y���E㬳-�:Ү�1�|0����Z>�Uw?��Z8j�cv0�=cl���={d����H'�V�{a������6 �ě�;x�§� yK&1�L/ ���u͊���+	Lk(���d��í �����(��i�D��wB�n�e8�8�şl �ey[�$��z��?-�>˘���ޱ�pd5��/�꾲�bGX����X���b4�u��n�W-�SE8_r�P�1�� ��Ȭk_r��s,�q�/L:�ł;�e�g_�k��*�Y�Hx|�c�ZǼ���4g����A�p�%��z��aV3 �	�w�m��e���� ����H�F�?�^n��V�hT�v�:ie�Y�Bz�(Ĵ��υ���C8G'��U���4�!J|s�v$/'��@��{�#PI-�cY�K��_Y�Ѱ%� +��q������Q\ܙ�����������9�}��x +Lp������45K��v���+��(���X_����:�Uj�������//^\�t����n���������0%���/^<t��I8�:��[�n���ė�Pi3b�������t���*)�C����V�&�OO��板�Ɠ��bRl�6���菊�@���ʤf�-�\���ϗέ�:p ��	EUU��TGP�P�������x��� >/��)c���9���ʍx?�詩��1:�&��#㬌u�ڹ;�T�d�P��a$3�WٛK��ְ��61�=��T(��LV�}�bb��[��ܠ���FTG�L�����̋���|}�⫽ȕ�gÁ������ʕ+�
,�lM�z$�7hK����`,�d�٢4�\в>N�N��ok�P�J}h�Z��W�o1lαjU���W��j5a��v�K��b�Z��f=0�Nx��=�N0^\���$��$�����i9j���f�J�a}@���2�I�b�F
�Cf
�v�-i�?|�fY��WF;��f/�f��\�P�c T�O��F*�΀�
�R������^3���r>�X�ز��V�T?�D�b$��h��uj��oO����혽�a�X���������?pӳB�8�ܔ�c����o���73e.��Xu��;��ha�(�J��J�<��c�\: ��ɇb�1 d�ҹ�X�Z��+o����	�vO@99���M\O�t�]���"�� [>ޕG�Aj6��S������u��d:��R
{��S��FlV>��Sc]����C7s8�JJ��=��l�����/�Ѳ�=e����W@�I�������4�^���jڇ�9���Ҧ�W	��2�4�b/�Մ�H�4u�I�`5|3�_�p���7da��t(�w>��AQ�����3��$���ua���9m�a��_���� s[���Ç�x�3@sOonH�NI[�.�a 1�u]��8v��=^���r���c�D�j��^b;?b��h,&f���ӪA\yⶕS&}%���c����7��~j��](�i߷�p�8�"% ]M��'Жe�1��Lc]G�&��F�sQS�}�M�6�(ޫ��X}|ԅ'�|x���X���J���c8�	�]�^K��$��de�	����I���~��t��"�����S������ˀ  �������8�O��?��d_��/_�����숯�}h�p��%�k�f)�<����q\ȫ =0��4l���r�5ji9��E���V�@g�G��0��!4����7h8���	 %�~���������{n:��B��T�������_m�]8�tn��pb�)�p�Z��P�!b�f�YM[��"M�ڸ���7x��^�LP��2oP%����@���*PD��  G����{�n/�g���W��U�~Y7{
��{�}fSA
�
��A��<���G	���<��)rU��?�����I�!lP����|3��^&l��J�L�]+��Ux7�RI������N���c�t�<"�[�S
��������t~�3/�[̱THtf��Ns�l�����3�GF�&&&�Jƞb�k�(�,�Xq��pD���F���<�k@�prAL��s�f�B4�};�w��`?�F�Hl����J:�M���,8Б�wU�_�8;`\Q1�v�;n���u��IZ�4��'r01�m�S���#�}��Ch.ONN����=����b0@��?�Np��t@�9>c�Wr����d��m���=��d����`�1`kJY�Ң�����FV�_�~#������yNNN����*�xH��߮�.�&��������˺�u��3������]�@�a�J.!�趄�(�&���uf8��h�#Ť���Ԇ.)WW��7�|��s�r���~tXB@a��O���h�7�}{mP�]U|�cD��w�` ��e�e_^�ExL�A�ޖ}�L����Ͷ�(�w����Q���1$y
����jar���tx[0K�F��[`$��"$�Kppc3�����Ev����oo�,��L���h*��QN�6��Ƥ�q�,�3�6a58�L��D(33�W�7��s�F�ퟓ�g�bi�
���E�XM�\� ��UT(a� ��<�x�K�����1��r���W���#̡�*�����J_	 ����e8�����	h8�f8��^qD�)8bA�Z�Tl���}�oX�zX����:�Q��u��{��.��ŞӖ]%���T�P�����U���N�:3�i�^!!2��s�@�?�����q�椾HM�D�B���`j˼M��@,P��5���h�(#���o�+(��$^ڰq#��S�2�������
Ԟ|���$�ùNV���M�0�Y�na{t�{b��8M�[��L���x�NcՑ1¹��,X4�?�g'�|�4���A2�_�+�	�)�����`݋q��ym���kx��֩�m8 R���Uǥ���<9tK�׭[��g�Ks ��X����	� kDXx�`3n�ԔK�n�F�b��@&$c/����$)�ceZk�7�	�BA&�O�P�ЇQ11�`q��}���mk���]��o- �S���K`�P� 2�=.ˈ\�$/�l:�[-1�U�Ra��q��>�@8"�Y�:]n]��g [�I�28~���x��6	bL��ΐj�q9�z0�x[3Т�H�}�N�e=�q%����Mr��x|��X��<�(�ݻ�Q��2<m���vefXNs~^�V/��ӓ�E]v�o��f�J�����@���oim���s�jg���uhY��H�
ذaY'�s��|�9�(n��zNNi����m����7���:���g<00[y�Ʀ�+����N�~������1Bby��X�uviϩg#����j�Bil��%����CѨ<Ģ���x)OsK�R�0MNJ����4X�ߞLăP0����í��C-�h�0��<���$x�+�݇�O|����^%,�����Vv�=<??NO/k2�zl����2��S�K�_d_'��Lo~����Me�5
4:�5+n�N��#���~���p�Ԕ�㝝��VV!M��Yc�s����>󅘮ll<��6��FO��Y��N��85�p���6S����j��`OCL�p8�afk�]ᧅ���|��1�9� ��I�u�
g������SB0�iP=�I�g�4���	����4��������R��f���"<l9�����oKqB�G�Q�iۏ������%=�Y5a{��UjzY ��N��$#C�Vj��)X�8�����W����n�~{2^�ڈ�r��pYz�I��:��y؝���2a-Q{������I�N�M��P��s�?�r��j��qS'��<	*����<�d��w� 'B�Z��J���8}��oLj�n�r���8Pyx��6���>"�4�W�"p��`�yxx\yt��3`���.2�����~����:w�X���"p�^���	���É�(�I}��*��e�8t��zx� ٱ�3�/'r�R�� `�\�N;ĠB �e�H�}�ѯ���������˧h���g�N@�������f��L_oc�.����������&{~vZE΁���Kغ��A�����X���ـ���P����v}�!nt�m ɧ�w�6�T��{^d�=ëh�����&�P}��ҧN��`�g������{���S��V�xA"��)%��w��1nܰ�\IM��"lD*FΓmJ��?em������A h����U"���,�LB��@�T ���g�}���,-aO��,�~E/1�+h�6(I;���%���'}��r�����TU-���1f3�����u��饥��$�ٻ7��t���ɴ�� �q5#}{�gFҮm���e v�m����ګ�}2Io��a�����7�]��0��X��>y��$�8w�\�ׯd���a��) 1��V>>>�;�&E�l;�0� <]�����twowͣd��F��.0&k�E|�i��49ܪ�C�������۴�B�����>I�����4:�ޟȍ��&p`������S�����}�
��-�6d��b�ap�2��a0R�{'gfܙ~b1��Oj�#_��,/���`xu�v����F
����FD�قe�-+Rq�6�	���ojj�7M�E��_~sx>f�u9r_���18o�SL�x{��^���)�WP(3����N��������)<��-!�ֵ����A�o���O�K#�v���Ko)e�>�d���6�Yr��XͫWi�}%��5�{���$�46|�va��������U�5˗��J�y�f�\1�3�
3��59�R��L*��UuO5$!�Z� �Ccc]�=�:j��¸koŪ��J�K�L�9���0���#�7��T򯚚����S9�~�z�I8`',s��L, "M�v�������L|�L8�h��ʥ}\X_bjzV<׳��_���V�:�t�(�͕,�r�g�����,��:���|��j�K%u�������xm	(s�����Ite��M���9�#���Z���@�:¹%E9]=�W��]|c�����+��-���/!1N��K��*s^�|�&["v&��7�j$󜾾NB���܍�8��{�>��"���B�;H�5S({�N���}|�#�r����������ǀ�����#��'ɡ�`k������&�G���g��1]5����y�R��e����8�lL���������&lY^]�ﾨ���G��7@	�sFWWJ]����Y�V0ܰ36TB�#�Y\lP���U]92��ee��~�@S������?���hL�I6z�xb�
c�13�n��U�Z�/ p��5�qԆ���z��H�]$VݯZ%��\��_*� 8NmY�u������j}�����*HNV�ԥ;�Q���Y�o��0<���p��~G�as���B�n��	�]!m�7 ��T����������F�a�J���⢴օ�a0���<a���L���)������]��(T�8p�������׽d���Zߜ��%���X�CS�}̛|��E��'�Oq	�ҮҌ#1��U_o"���᭱}���,�Y�96�9� �*��N�J޲�f:�P�V��FL�~H����{��Κ�}��1N���G@<�t77�]Lmb.A�:����u���q��)��W�U�_�L��\[RԱKޅ/�$6V6�hq��Ag�������њa�u`��b6r�j��'@��?+0) �}?г�߇f9��Ԣ��v�]Ȳ���������7��x���W��08��.߮ϽS 6#�����m���i��>���w���,4_ߠ4��h��ٳ�����ş�m.��W�~��ޟ���(��P����+w�Q;\���һY*8�u�d�-b9�s�}��;V͗N����v�s�k��O-��x�ɷ�B��g��ݯ��w��?���y_e��=���/go>�s�j��[�{��*�޶��]-SM����O-d8�+�,e�#֐b���#j��3�\��q�ٵ�]��z�5%�6a�(cT}��}��g�Ai�"_^��WϡI�dm�{�Ԟ�������<
>�LUW3r~�+46 ;_q���ÚH�M�<��/�8Kz�F�C1z�WXx�\�ڦS�wpS���|�<�+G�t���P�Ty�w [��/�ܿ�x�0��UvU$/�}8Fe�Xg�A'��Ҩ�E���Z���ڶ�6�P_�zS����-��=[wp�������4*��遦��?�]sJ�+`�z���ʬ�������p-`�mD�χ�t��7G�N��돸�6�J'�&�f��c��w/=_tlM�K��o��� |���Qt�f=���Va�R[ʖ�b߂�R�Թ3�r�ڗ׾U/.�)��$'Y��IK �ô�-�ݍ7O�]e`�~4�{\
���l�f_�*��OF�o�-�}�Y&�+��J�=��ݍ�h�4L-��D/��d?��%�p�z�n,$�фC�0<W�A�����[a���Ǐ��+%�D4�GV{<
��J�kʝ�%���|��4Q�s(����c�|CE�cc��'��^c�
ѽ�t?G�E���^��ވ�K��3c�Kﴫ�M�pf��������vr�}�STf>/QqR�WKmʓڄh!Le�L���Ɇ�Jl6j�{��E���U�L)�R��@W�o�+���5�6,=LU�{�yg#��@��?�Bl��C�/�I�0/��;�Sj'c*�Y���;�	(�>��}3J�J�C0�e&�!L��+��P5g|����qW��T�e5H���oq����{�s�Q�.־8N��ǃcx��|�~�Ca�YO�	����V�5n�rc�D�U�|� �]4���8������8��s�Fip����b㖴��̴�ISI2�11����A���I_�0�y�M�s�QV&��X�-�����.y�#�w�4<)@�<�wz��>g���j��|;%����l�ف��>׳6��aУG�Q�����4y#������?T��|�#a*�p&���궫���W�������D���k���J"�!Dϐ5T������48�w ��-&��8+�M���5K_#�h��߱�~yE?�2u��l,t�V�b��q�1g�B���?2Ϸ�f���k�}�7?�m{����&C���!���r�A|���=�7W@)�ᝦ��k��>�HL0�>�q����4�r���2�،+]=%��G\(�wO��^�x�VX�ص%�ھn-�̂q&?{������*[�����jP]�C6Ol!o@�_~�Sr^�xܔ�AN� ���'E듹5�����������c�2G&��@�v1HC�Y!X"#iZ*�:�����m��4�
�⫝̸S��k�7�}�q���899����q�&�� �a*�	�_�&���0\!���)�xA�!��I>#3"|LP�`C�܋�(����:D[3"��M���~��SU'�N���׸�PEi��֔�-�\��L�����hZ|�Yfo�D�{؋0����V^]�@�5�	�<�����M��x�?��̦�c����3��Z�YU�45�#	�Y��GG�?o���&;�_�`����	����t����S�a����G���H�B��_�|N6C��L��:;�{�b����H��E��+��(x�;�n��l�vbc�Z�/ �S�ٹ���G[BA�a�8@�f�v+WM{�\:�40P��&q�,��ߖ�}��ӥ�!�=���MSa�0�Z1R8=;՜�M&-v�9Ĥ��m �W�&�.�:4�6Z�)�|��k��ȧ&H�?D��5�Ņmބ�� ϓ�-l�P�?�,��3�_��۰}g�][�)��eGD����E�*Ū?�|�6}⹌��B�7�6�M��
Gh��|��@��Ŵ�F�����i����N��W�:�9PߨR��]]u1o8;[��$���2� ���$7+{j���N=�Df��`�]C����Sm�X�����칏�<|�쥤��Eˆ�-x�Ex��W����ܴۍ�z'�k����ʔ9p�� n��A�i��V2�~Q��.���+o��+%\��`�_�{y����k'd�Ǳ�ħ������_��}��"Y� {�?VL����9�	H2��c��V0P����#����p̈́,`����wl��DϤ�\Ӂ�ؕ��ש����W
>+�\\,��b^x[�'߹J�H��ťs�"X�<���v�c��mV�L~m=��ڭ�d��ʮ���Ӵ��C�@u2[�s���u/�h-2#4#���H;E}��|f��-�&i��A�_Mr���,p��3
��*���Z��dv�*Y��_7����U�*IO����T���%h��(֟j%��y�r8�-�`��AJJI��0�G4� 3%����l��+O���b�)we:N��pD�r_ǽ/tyO#c,��>8�(���2d�J��&.�̦�oo��^��IJggK�XIz`�*�U��y���s�kj  ��{��5 m�^���@vF�ak_����x���&44�lc�)���}bf�,W`��Ya��`k��8P/]��U����*ց:�#��<���vU�r�㧹���G&��[�<�0�ݴ��u�C�fBt=���m??軑#��:��I�i��zq�Z0�O��E-�w�`0�Al�cW[[��� W�bSGG�z���̄_�����D����S틏������P�V�����e�n��i�<�t�v �m�g�ToI�!G6���^�C~׊����W���������Z`#�	�`�}��ؓ��6��d�Η`���mbS�y�ى�]޺��\ԁGL���O�<){Z�XT��d@۰�� 0Ʃ�\�~`���YJFt��εI�P�<ODr]/�H��e2��j��Q���+H��zSs�R��j���,�U��4���#dSAW��.v׃�UNH>!���������0��9�r3za��� ��}Q: �h�B�N�`������������j
T����/�kÅ�a*��/�������Q�����f����p�ƍ�Z?�U���DsB�lk&n/����C�F�8��E���[�Mj?Q��k��b��'�F��>��!V��L���n;�7�G�%�o,�N�$?V±�t��JƜ��5	U�Y�<�0{�D%��K��1�� ~Ԋ�J�^e�922873q��k� tN�Hy^>��U��h��Vn|
�%V�P�{c1\�Fþ<9��UH���܀�kf��d���R%��wQ�|�� ۯ���Q�^|ףY�8?��?�J'j�:�/b!y`c��/')]$V}�9f D�Ш*v����>���<6�6�����u�6B$��6��;�/��TN�O���s^�:���v
�ޢ�݆�[�zT�����W�sδ�G٫˼���Z^5oę�q��&\OIc�������~�-M��Aü��[��-%6���}����N��¸-�Ί���	��#J��ٗ�� ���yĥ�6o�y,�̽��tD�a����i��q]i�+lR�ڽC-�𵙪�ݻy��J��3P��g�<�V���Eq#��PS$-�i	r�~�,�Aɝ��;
��2B�S0��܀���3;�ݿ-{���	h�e����I츇�*�<�ب�G�=*ր	L�\}Ȱ����
�k0��XoA(	nr~���� -�)�8���皸Yc�|��
dv;�@1�m^�A�Q\!@�^�ų`��l;Dc�s������k<J�&��N��߳�ټy�e�9�Hlj����8�-��<R2�g��%|+|��}$w���;�̻�6G�T;3�5e�����u&�nzw�
�Ye�> ʬ���[��X�\ug�g����/0�=��3Z�ֿ� JgÓ�o/ю^���/C�KU^�������Z*Z��ښ��P����^7e릟f�����1u|��& ��vk��t�5>��5ES�Ǐ�D8h?S=��=q���@@��&�s��a���@%��u̒2'��d ����V��������ϟ��;�~��F�]��P�f�O�����ߒL����e}����k�h�̫�� �Rd-��[�0��^l3�`]��҅��A@��Z���g�K��b�-��bM1瑞�G�����ڲ8W��9��M4��rν� ��hdH��\k��c��c�n�+���6�s
�}X:3�h�ͽ��Ft�|������Nv�,iz�E�@,�Z�*%�)Ϭ<{��^��w|e���/����%��L�Nƙ�gv���Fqxx�j2}.�b�τw��%���O��Fb��{ ����9f����6NF�Ε;3U\�����-"�3'�BG�p]5e�Ҿ(8�μۡ���:���"CڈC�
��-S_�
SI��?j����x�}be^%v���G3Ֆ�q8�1|�oZIs[���8s>��)J�8�n�Ag�{��-�67.oU:?b�������N�,��ܶt-LI5�����4�&i�SNU���������s�t^��B�d��/�jb��<��� ���?~��uQf�8�&��6E���E���i���+��w���oH�k������d�Gu�2�����C���o��2�y/���]��~��K�������
o�w��]�������$��s�[ķ�ק�;�_�q�����cTnFU�@V#hp��b�hp>�0A�V��t^������7�b7�@��4>aD�t"�o��nfb��!���u��N�.���:��Hu� ]ح �!� q[f�<��D�T�Ⱦ�k��)Xy�KC0L'ׂo{��[sB��5x��)f�bC쯤��΃�L1��L#F�իͲe��qM\����^��a�4v@��#ܕ�����v��65�P���B�:�q��۩���d'��z�H`�n+��.�_1�)隞�tR�(������i����O�?.p����Ep��aE0x���z3��22��	-'։�T�g�}}TL��&G�fF��dٜ����ZcL�&ڄ�5��U���;��S����r�6��cָ9���grc$�w�oZnbN�{�x��hru�ui����pp��9���.���=���@ΰ#N,�����4M��
6e�����婪|�se	��>����Ql0
j�+*Fʊ/NT����m���=��PT$�X�S |1ȏҨ���f�3�����[��^_~�y����Ba*;����i��l���ɇ`!��JFc�>���趭�xRu���0��,�8�?VI�]O[������'�y�g�`g��;�F�����+�88C�w�4Ps��'���'�/i�ħ ��=Xe���Z��t5f,A����G.�����v�6Z���.�N�e�12�g'DO��;��4`v���`X�D�޳���!pѹ6�te��J��3�(�e=��LײrJx�e�d�:*���yx����|Ɓ\Ƕ�%�m�*޿�i�K�U��i5~F���9ש�?�u��+��̴G\��8��N�[�S�"SGy{�����/e��p�~4����|ላ'k�w|p�c���G<l��#r>�~ȡ<��7:3��D[(��D��cCav.UG����8�l���cN���_���t@���^��B��_�_uR��5:����&�u��B�_N�m�^����X@�u�ڵ(�}����_��p�����PD�|��eOgf�����sϊ�(�����i��E���{�^&��8`s5� ��u��6�T�`�܎�NN�4��	��:b�^e�`D-hU�P3�w��W���ͽ���ʼ
�-UIz���+�d��W�|�ץ��k��&�ʮ���%Yi�A��|��#0{�p�ހk:R�IF�Pʁ ��]'��1r���9ZY��6vv�?�K�2�`��!�L2:b���uV��`�w��	�+L����#�����9Y����*+�	��}�X��V���2��,��Ӵ7�%mS���Xt
{,O�)Nu�؀rc98�Q�G̮�>�zg��Z�ѭ���q��n��v�S�W7Ug���~@��]�l��om%3g3����y�S�
�Mf�hcK���;J�@6��Bz>hz�!`X�>֠�k��L	�$1�]nq�2[90m�HD걶��xu�n�Z�>2S��%eU(75:��/z�	����<	�8�����/b97[�� K8(j�y}\@���Ɔ�g��/���5��-��5��=\rC�Z�`�g��M�>�ǵ��l�h ������rOD�R�$Kq�Q|�	�Oǜ�b�t����|
�wj��ĲR����~\�ǅ�cV5�ʻB��P��L�� se�u�'�p��l��D�Ϲ\+Xp����Ub���0�<�v�?�yLά n�QZn��p����G�m�á��~���f��gY o�i�a|b�	�`P{����V�P3��5Q����'��]|@]�I8�ս@� �ꋔ�ݦ���L��oP8���� ��;1س�3��Y[�a���P�q��ۈ��q w��x�x���B��
�������BR~?!�&���K�j�=E[f��5��O��	���}U1����.�� ����m|��qVU�;Q&N��õ��jM�[ɘ��.����d��"��U���bh�?1���XG�=o��T'�h�9�L������j���J���`�'������,Swр�3�Hg!�5��{��O|�qr빹��u�9?퍬'v�����ܞ`es��Lx����/��kX���"�Ƕ�LT�8��)�x��_e�M�!�0�6"�a\�\������ d���|?��_�,,d�AT4I񛸺�"n�P �⏂��c_��]0�!W<��3���@�ɓ'([�^t�pP[G������W����s���a�~��)����q���6�G��E9Y�\��b���=�R���gtuW����1ȸVc��B�����P��酫$���D} ��2�$��d�v�Y���m�*;ؓ����c�v3�M��>N�ឞ��[8A�_��@b`eeu�w&3r(#G�u�p�>f��#z�ňnE4VDt��̔��:�}�T�Ne�o٠u 6�#�_~��m�~�r�9�xI�8 �koh�6����S�wa��h �'�>��9�L.�� �s��^�ǫ)��<6�S\l#c:�(�ѽ��q�I�e�)B���|�l?�x��'�T�=A~��{�%�"���L��������E��~\ ~g����}S;��
M�� M��&�Y���YJD��U��k��N��\ C����Tp�}�k�&�̀�.�6sxm�k0H0����<5�0��k�{�wn�$�[��!g��Jz�'#Q,)7��*?���5��@Р�ܤ��䲯_㰑'�j�-eU�5��gf�Xt���-[�ǿ1���N��.@��؜%t�ʴRCKf�V�>�tB��f��H+��s��������7�)��P�c�lc��3%D�8���/yEE�J�	@'̲S��v��v/9���ͻ�<~��-E���R�FGFA�L��;�휡��>/�YKA��Bf( orm���X�'ݱ�`_u(� ��|��U_����Y�?WtK�Ƃ� ���l������+�7�����Y�.�M���M����Z���ٳ� x����_-$�D��;DL��3R����L�-�NNN.o�{�6�g5��P�$��0c���_���	�:�v&�����z�U��V�0�$�c0���d�_eg'�f�IO2˞��͸�-V"���69����n���w<��v>o�n`
x9/uG1�v��@��]g��i�_5�#;�G��ݻw�n������'�����m]��"ķ��������Ɣ�p ��"���a*��}q�ao�\�WHHyv�r@Fص�ij�d�j���&==����g�Rb֢{vR�pj���$ЃN[]ໂ�<{�����E�L�Ι�R:]ϙ���R��mr�<�1j�ѕ�49׌�;L�*��N����1�`���A���;nYҲD���u3����qr"p���}�c���!e'�.��2���|L��&|r9�mּw_��J�1^�N$7��T�U��q����*�(��Ȉ��y*� �œ�T���-��T��T�	�E��bw�_���!R&}z��_=���055uė�zfu��"@��P*�o�yQ�c�� ��pA�ʄ ���oV�M�|둭.��a"����li�r�s� �^�����p_�7v���Uf�p<��܉��C��ɱj�].R�#��+�Vf"�=D���	ZbX8S'�xnL?ޛ"�
DC���_�}؞��酞�8�x�C���h��l�mW�\�!�u��2�w��r3�R߫��I�_��d�D?^1@�p¡2|4�>.��\�U����q�SL���v!�o����n'�� ����杣�Ȑ���1�r׼����OK?��Lo�D���B���ʀ8�ax�,�m���[��)aaaew��k���B�pҧ�	-� ��s���_%�{�9��A`�1n�ও�+]30�(LhK�t��坿�b��+g�I�j	��)�z�������T�L�jb�Q���~�6gL�;��z�{�ׄ�+[��	b�� R��8�Ⱥ+��GǰX�� 5`������8���p6��O��;��6��i����9���wq"��C�jg%2y���;��2k�XdH뗝Rk���;��"�a��ڌ)K��۩e��J�����劊[�1G"�w���'1oc��0f�fƙZx������\��*5�|3[s���e��z���Q��F-V�0���l���!)U��K
t�r������b�#�v��U1��1�z��e(��b,Á�}�>*��C��E��pl
db���с"�#�<GF�+�x���ȷ4�Dl�om���LV���Z��
G���12�1O;p?8���p&�n:�lL�]��`�6܋a�{J�:b�k��D�86�g�Z��d*��GL�l+{�&�"�F��۳ ����ka/-+�g�껨��Gɿ�����ppN���&d���<=�n*J4̌V�T�^�n��(77W�?�X�!�T���8�u6�	;A0>.<G֍K�^#��������֠��W�l�vzˣ�S.�
>��y~E�����ߗrLYY���BB��P����'Z
�����+�1Z�� ��0ƭ��W
��msmj'd���I׮u�G��k5���^sP��^����V_�*7>�]5���J�k#r��Md��E�t8��kXd_nX�8��r� i�@e���ڹ���^�Η�4
�����%Y�c8����"�`[�p���8N�k��J�Q����c�Nj��<~ٔ�%J��AO�k�Y���s{j�}�!���Y�pQ'�r�S��nƙ���M]TL\�y����-�J�xX%q��Qtt��e�,���]g)�iab����[�G\�E5&�h�-1�"�����KCZ�HT�3[� �h�Ӣ��4�+_����BfO�Q�ҌöΎ{]d�<��5c!o�!L�� �p��/�8����87��
KC�h�;�rR��F��,e�'�xȓ���d�]jX���(�ӏ8y��_f1A���������JF��/2��E�q��H��M̈́��C��6��q�#����n��y铓X6�F%P�$�i��+��N-����r�����	��bþ��1��*��?��,�I�#���H��MGG��F���-���t`�� ��Ϻj�@��,�F1�̽&g���x�R4�?�ٲ�W���!R8�: �����I���$ HR��(S��� `R��唦%�2X�m�M$\祬�a�q�7��2
Xdxp���wf��[�>��}���Jbp�DMv����r[�jl�U��i?�K����Noa���)���xdý�?��~To_7����� ;���7����{�M�����>�N���,g^P�А��}�U?�`_�	 ��7������D�O�I���^�4A�VG�Pf�|��M
�QXPp �G��H<���t�-��c�ݜXc�s������lP|9��(��?a�AN�0CQ����{P?�E���f|c+@�U��@�惞�~��׎O�>鑉^�]N|�?=8=ee��8���F�5���2�h��1<�me�J��`KC^S>F�/b"�)G~���-1��L%c�Tv�0/���#���0A�h
�I2����BD�Èѧ
��W��ݞ�}��0��n-�>��֒i�hz������(:P{��`*�}\x%@��y1@1`�w�x��I����X<N^�c^Q�S{藷s�~�"�.�>V��]��q`yj.� ��'Bq�W�@h���Dc�����C�d�j��	��7��?��E�'���J�&�g��=^�;�X����t7���o<x��u�Ә��3���l�鏈:�o�WC��|�d��싽J��pA7�	yb�3[�A�\�v����_�����l���[�}�֚?~4�l���M֭�]W�,S��%�m)ǽrޙ1iLr�7����[���k' �F���[�00D�n��$�42!�~��j�R�-�B��\��-ͦ��L��"�(�<Y���\��O���͆������T�'n J]QH�_��i*�z�x\#�hc����o^
-�c��)�0�2պ=i�ҤU��됪�xT&�^� ����*�x��b6�7"@�n*��\�9h_�A�&7���=��{�A�����$������J���4�k<���f����鮶�|�6��}Q8��C7���ϟ�I� �$צ�����ӧ�R��F
��-��;��Bb��$+l�fy�6�c*�	$��h)��B��}��U{�-�B���b8z�M˙�.���j���"h1�l�g�����~4ݥ5 _�Y~������%�I	WIr�+M	���S�@�A��4�}�d hԊ����B����f�g���,|5�?G\�,c�0����q��T �I���"�A�A�Ȓ:ѝ�"n%i=�6(������Ů�=5=l�/�zgz��!.t��7M�<G��}̧�F���E����d�� E�u����5��gJDh	�q}�l��:�܍,�K��͆eW�FgK��!�� �J�l�/I�|0����'����8X�S��U7����������M�DٟoE�x��q)��E�c�ԣd�=K�vtsx��"��"!���7���|�`؊���a	$�p�c@��֔ϩ�)n�����t�A��I7��fm���5�_�������@ã*RC��!��|��{����9��Asg�+yQ�@��뢥���������s,��5JG�2N9���O��Ϟ?ߔq>��x����^Q�G��P>?� b}>�9J=��0�F�D��%c���]��X���"Y��.Q�@���N���f}��z4sΩ!��@n��$��ө:�ݷ�;mu1��GT�K��N��4� �㬪��ueeގn���vw�M�t4\ފ��s+���I��\�c����k.{�"C�5��bW:�a��>�_Pӵ��-��$x�����^JR�&����h��w�[��m_���,l�~k�ui��mZ�"4��s�Xx��'��:�.��k��n�Wt�v��T�47 �����P��5����� ���k�zQ\@F���'*^�<a���%������Z��T��Z%|[��ӑ�������S����í�r�x؏��+�s���5H�yhC��G�-���-w˟��H_�w��o��N5��k�'�z�2!���*Ĺ���-��wh��S9�sn鬒W6޲���E�/����]� �C����?B]������D`��c�b�&�#f��3KCkzN_�J6
$ؾv`�C�ހ���X��c��u&=as�4�{��RX���ax�+'��ƀQ�Bi���o�;���K���dB��m0�=+z�Q����V�ڬ� �=x� �-7 ��j��5%���O���?��VJ���0�2�����L�7�	?����fk�kI���C�N��)���D.��oA2�;>��.Eu'>�+kuۗ���SP����������2�)��ͽdUM ��c���HD ʠߺ
�+F�zo�����=�s"��? ���t��x#�oZUѺN��FUK��9��_���@�}��~B��hű)<�Ct.���� ��e$��[`��s�<@��'3}�v$5]>-���c�3A�|v�o���l��]+�1���X�x�a����Ʊw��c��a�i����W�jMi�
K�#�#f}��lXx�T�Fн�}T9��\}Ȁ;�Ui��VVVC�28�:ҥ(�0����wm>�{��Y��]!X� ֒$ibY6�����
����%N���WG���� pu\�lm��^n�/�T/��ŵ[�/��+c����|N�xw%;��Bw��HTxbι���&�G<��%x;�pq'-эT�O����^S_�t-Ey�1����w�۶G�u_+����\y m_�~����ݼA����O��"}��-�R�t�7-/[4S��Ȍ��-����M��d��Q������*�Lޓ�:*5����G�E⃣;6(�7*��*w�7��~�2����s2)z�w��+F�.�.���2g������.E<�Jۯ0}5 ����~W���!��÷�����Z��NO(#���"�'�@���U�?np.���F�a8��K_����ʵ{�7�$�Eѩ�v(c�S�D(EeH(e˴�9C�Ŧ��$d���HR�v$�I�L����9���?���{�gXõ�k�{�7H/�u22�P��p�ii��X�Ϊ[í>��]v>b��W��� �g��H�����v���/Y��q�������!!�N~�t��a#�0�Xm3�MaeP��Baڍ�V�a�8#�{\9�w{����np}�������qr�#���&
�U���>,�HГ~��b�dF�K�'� ������Ԛ;{څ-?�~��Y��a1���kдFߎ����z�7�Ed(c��%-U)������^G�K�ːO�Mw˃D��`jm���_[B�!e�eCJCT�D� }�>��Ӟ�����{��$��Bb|���n �;	&�:�fGZ�>��L�������kfrj�e��@��{vƝ�ȧ�<&D�kX�~��M�V�B�Ⱦ��5���'n*�P�Kv
= D"Լ�)s�Z�GD�Jҳ>��^Mp�\/�[�������#�a]���mcS��b�5w­��м��Ua-� j���^]���s����4"}������û���{/6;�KHĖK_�3���@�8��� 	um���qa|�	���PPfj��[T�9?4��֦1�u��X��[�$��d�Ic�n�3���k�g-e͹��a��lӢ �ʥy*��=/�`|��@y�(� �z4�>��� �I߄���og�:��5/�IF�kf���2U����Kwٶ���lc���1�͖�L�]���O�Z��/�Xm]��c� 	]��j�A������5w�L8�����i_��p��eAv�"g��Q���5�pc^��-[λi��2����C�V���?�|f�;���Ç�dggC!��u(����x=�� M����B����N��Ȝ������?�`����o+G	� ����N����m�%ZI`�O��F	��ڴgτ��R��Zb��=�m�gK�p{|R��+�_>"��O1{�t��|���!e��T���h�`�z��m��n��D�uꏁs[���=h��o&�2|K\�(/o�OʹVRR2�g.�}���W��KvDкx���:-B�b��� �G�Mk"׌��/[���)��Ӹv�Ės�`�I��a�;4��m��l�P�L��Z���G�&��عsgNO����---��%���Kcm��k��J��1�u�=o;4�#����x^r3��#�ի{������7��vFܦ�Z�� ���kmnoWb��(G#�B,���j�׀0�h}��HS�N�������iF���D6��3�mt,)���m�aĹ������� ��@�x�L E0�]�5�T	r縙�r�d)u�BNu�]��ג���1��Dn��Apn7FOkp�����?*�26\�S1na����z۝)��p) u�d��)��X� ,��
��>�"Y�P/c�����d��NM/:<!�\���A$'ge�⏭<�fb�[~I��եW�l2{	�,Z���gh���,����I�M|�]�V���B��S���/_���3�\]%g��.�s�{.����c�
��wC��_S!�N�;�� *h�iˇ�k<��R���qgO4DQ�X���qa��xcQsQЂK6N1�.�ж�sw�|�2����M�Nö��� �aW��:$hq�G%4S����`�b4� گs��YYȂL�����wA�#�3��N�_`��H ���%?7�
4������06�aQ�������,�QKOzN�6 o/s��vPss3���[RC�{
�-��s #@�]Ќ��v�Z qS[�En=�X�o������]��3��]|��g,h�d�ç���n&7��]���$�P��H����~H��2���j�IIٝ�+bӹYe��INIY �@j���7dʇՄ^�P5|�8�s1���\�;�0��I���.�_�4Z��*�v�@%�~��E��l4�,����JK����[ƞ;\����vQQQ��O����+�Tv�b�&	x);;Eq�n�H��f�	)x�������d��A��o��dPFN��q6ْ;�����\��޶��6�w�H� �GS=<��\�J�50����1�q2��`�fV��~�`��.a��S�<�F�������E�w"��p�Y������^��h96������wF���M���]2��=�l�5\T��M3���3ۻ���d��x�:�qG��M0з*͆R�L3�\��Um���9.���4�U[��i�����s8wn�d��D����^4�6�4�	nw�	�� �	�U#}Zܬ��!%ə�b��ि �(,�k��k����g��E1�a�gu��n()������xK*�ugΞ=��:Uϊ����7�*����劵�Uk7/j���i���3W][o/So����c�w��i�� �ߌc��=�֯__��`�nݺG�f����pV�I����BM�5�KL�b��|����D�_s��&W��8\3�r<,'�Ѧa�&&�{�!�a�m���P���(��{Lq��緎��g8�>X|y��!��Ûc�^��ؚ��z4֐� o_�N��rSm��C��k���X��������
�Wq���TpR�Hh!��	%-n�l�o�h�o6aF}�-}!%%�H�c�)/��e�ꞪG��p7�1r_��X}����!���߿�����Z.|S �����=l]�͠�M���u�&�S��̥2��Dx��CJ���}:E\����'j}���k\��i/^�s]
�T������q�cm��pJO��p�2� Kc�PF�XYz�^�#H�mH�C�0EsG�rn."�������R45qs��p��)%1E��ͷ�W_Cw�8�է�%�J�̧Sײ����Y��~��Ձ@	�������.S�A�f��3�J)������!P���հ��*�.�7<�q�ŏ9���*� �Lt.�%��G��Pk�mdF��r�g-����̙3�� ���5=���*� ��DL<�:K�n��7��홪�!!!����+jAL ��<�Y~��Hc�=�X^�����A򺒇@������H��0�C�����wK|ƹ�mwF�ϩ�.[	�K�e��+6���u�����+��㇍��0_�����\G�hx%��k��$ƥ�{�$��A���ݶ|
�U��Չ�BV(fT�\|D�q���D-��8�YyBBB���$�e����� ��fʓ �����qc�}�T�ۢ�7,.���)ݭǘ�M�w��9|��뱵���i��<>��B���1��,��\�7�=ll<8�S[��ߏA�#|��s^�Q�t��C(J�?�O<�
D���X�J5Nj�+��|G
Y#_\Բ^�i�֑B'N����~s�45=l�C3姀�h���ȱoR���v��2�0'�y:��!����vf��!��`�)֟�|��G}���~�~����O�ј�W��}�|��}���!��z£׭�Mo5��C ���Ռ|�[uu��`{��\,a���^��5�T�]�͉ �t� -�ɉ Z|���7U�:�V�t��<�v�J��2��]�M�+b�����8W���Ąc��1��ڲL�S4�`-B����^�#
6����ڙ�X��U��xM�\s�Ud��C���
�b�n����"�Bmt�f}��g<��B�mÿ� �H	��>1vX+DV�m<?K�4��ܞ����u�$%��#^cO�|�ߕAM|�þ#�g~?x.��o��w� �cF�VX@��V�]];�2�m=_���!�Ŏ:R���f�� ���
͛���2�ťe�#;�����ǒQ�Z�0��3�tT�r�=���:��R�Ha J�~y�hEd��"��=F6���(��MQU��T)4�X<->�U
�����4,,�v�*��.B�!=�9�/%r|�m��;�m�t�����@=)"�턦��"DŚ�h�=@1*9�����6Bu�j�t̸�:�v!����7��m�}��/!���e�}U4r8���ӧ]�����j	u�r��+�m�~y�}7=
��tmmm_U�<E�}��Bƿ�L��TɔY�kzg~�|�ШCOC6UĤo@��{7B�Z�b��<�̿<�����L0(9e���eK ��]ttw�6��r��j��,�h�!���Xϯ���8��:R��ы���,��>� N�k�� V�;!9G�'�$7�9��)����[R:�F�E�9��#���IE�q^%|X-�E�ݺms�aCzk�4�L4�4]V{�@*�\�"��opL;�{�F��3N]X2::j�^��6�q���
�TU� �JC4	+���@a-��c��mw��p7'���������iV.U�Je�'ߩ}t$J�>��9LyKu�N�=�t�����4���^:ƭ�6�kju{n`�j�Ԑ���n�������|Q���	��|�Ϟ	��_�dOѭ� Ħq?rrqY�_�B�����L��ǚH���+������U��,����R��Zr�_}����;��x��@,���� ���%��+*�~��=�������Z
//r�����f ��R�n���9�~��:�{Y��"T��`������G�6���H��X�"���U����q���W/ �l��>A]�����|������Gu8������5ʊ�[!;;;ݓ���`U1�M����A�y��nZQ���a	�S�����_�M��m�w������ఉ	TW����a��Bٗ�nv%҂�pS ����ṯ��3�߸$ �Fhұi�Bk�:��c���os��ں]��$*u�㨋2�}��A�#�H;��o��T <D'�tg��+�.F<O���n�s�s�+S&���Z~#>;ܦ����3r��V�' ����
̸�
p��)>�����n��5t�E��3Ra��8��߯ ����Lv߆Xʛ�-��g<f5����6��e�$�	�~�����x��m�m����a��L�E�&>��AU�WInȡ9o~���
~���� sL�	'�+�����F*{ǫ1���8N��`���	��|��W��ʋ/]/�qo�<$d%�wϾgllP�����rL��e_��ev�N�P�]E�� !���	�Am��"WѾ􅸪��dl�X���A
!��������H8�+�F�@�F6�lb�%)�ÀǥT�s�S�6��|_F��'�-���*G3J�X(�&,�{�9*1tx˔~4��J�)���Գ_���<�۔�x.{[L��HN��ۦ:��b]�C��ePQQINN��/��a:L����MM���KE*�.$�O��ym' ^�e/C2����@v�z�dgOO���z��W�S�䚯H9P|�B}R�T�HZE����5�)jkk��z�5������oZ%QTT���ń ����D+N;vAff�n|�^��	�E ��_��60շ��3�4��Zn���6Q���Kt������Q<A�K�F��%DvІ7C�!m,g��uć닻�d�r-�UZ���j|�k��㾙�#�[�j����r��Uby��}��m�t���ѣ� D(N!�ǄE]C�k}� �\["I��;�<���N.p��/-&�:��iBB��ml�a���@d�5Ե�1�C�C�N�>��bR�p$3I���rut�5ZP�⴪��,'g�4�`[�&ciH�R֬Hc��n�������o�t<W�&N`�����$��4�3�f5�}*٥��*�_!f9F�w�q�|��6����]�:����	�S�9++)�ɱ~ ��};�Ɉ���&�:`�(A�=_��_z.��V 4���l7���S�B�ܔ!΢!z�槻t y�n�f���R��Ȭ����?�'Z]QWmZvzс�T�w�WP������׹>��7�2�#|��0�����}���<f�zO��!*CQQ�A<��	L���|	]�,�+'�K���d>Q�kmm��Q�����۷�T�/2W(�����w4֜�LlH����?�kW����m��� FZB(�v��Y�E��<��zZ?R0�T��PY�H�k�fr�� p��y�ML7�~�U�Ӝ4ў�P/�Q9.@�V��~�E��v����n`˂�� ��؄����rʜ���]�<WB\$k9���ZipUU��@�AN��'ǌt�\
և�����?�#w�?r*�rϴ�hރ) �p��5�'O��3�����7��P��+��U]�����럿��B %e� �O�qV�����:���Hϟ�A�;,��hm���E+��T���=��J���Ս�H����)�1H5��&���/�m,31�;9�QT Ӵ�5k��6��71V+ G&QB�s��K	_�yM,k�G�z��Rx�(�KJ�I�_?tw�Nt`~���%��xA{��}VVVS}x,���۰!�	@��TX��m(�����!����|z��L&sx��$^�&o�Ӏg`��� �1��Z�Ȭny��U���G��y�����.W(;�9��x
rj*�0F����,<�H RM�R��� i���^�z�\����
�	K�|�T�4H�VK���@�`Ė䎕`�R�W���(�%)6T3�T<�.R�T9����-P���FSD��"=��3~�,>,+��	fj�X��| ��ٷ0>�5S]zݙڙ��9�&�� 9;�-�����*"���-SN��)"��r��u���ݝ(�H�`���hPE��C�8+} ��"!�nYQ"+cK�%,�ڇ��mVL�ϟϏ����EV�.����L��b���'!_Y3�=�QH�I�-(3�@k8CЬ1{㫯���Qp��Hx��H ��}�1��j�
}��N.W��#
'C�+�Ε��*��Ƀ5w��t�U�F6B
��@�/�3~l��ib�+�y����c� r&~�L�"�b�̉��b7pZM��ϕ�9�w9- ������SF"���� ���L9T��/`m3�E=v�	G0�4c�
�b�Q�,E�L��[NDA���"N3�9%8����8T�jG� Ғ�&����$�9��=�}�4)�Zt�q[�)8�Q��� �41L�`���I5Z���z��I�w�ڒ��j�����[��5�ҧ��8���]�YqA@�&��� �U:� %d����)>��7����8�"�T7 ��Ν;�2��r}�!�KU�v}G��  g�#6 d_��>�y�JY
�/Ϟ�P�6�	����F�5]j$ 5�鏘�p*�T1�Y�$�>��G�D�r2�C�(=��t�2j]NsK��n� �=miiAY�%C�W����n�6ց��Vs�`g��c{�u�80��� K%lvs���)o��4�>~��&
��>���TR�*n�� ⅅ����G}[���ϟ���+����P'$�?��:���!Q`�*"Rj{�Ɯ�2�&���.��7o���EM���*"�\�j/ZSS���c�>e�r��I�",r�ܥ�VVH��I�l[��3���c'�C��0_I�p�������J��g��]EL۩?�+(��IIIm���3���Tc��1���ٜӼiy��إLu��	�N@����.���R�_������9"J�^��h������k�������J��E� m[p��U��Ȍz��A�O��:!s���2k��g�	��i����/��@������I��ԚBQ14}R�����ܚ����=�#3��n�?~B-000���bb	 aG�w� �W���9�۰������8�sf=NF|��'NDP�˭�Q�D�8K����Π�_y��T*<.c��U������ ��^(�}�<?jYW�	���f:�%iD>�/<<��N�yT�搉;pn��>�����y�2��T06辒ńU�],���������~��m���=�`��d-��]�I�a�@�}��K1Kb ���O1��q �P��.ݽca謼���F�]�& ����=jl��I�9촖�rA]%�rN����@�}��'��3�-���vw���T�^mja�8��k�G���a�����zs{x	эU��Q�o|�i��Ῡ����۴}%���>_��E�Q%A�S�M�wW����*��V���A
U�^I����Gɮ����2�r��} {���^�=��!W���dV�\�4\�w��NZ��ZkE��i����K���n��B4���t�O�k��bAj]xr����o��Ð�PQ!�{�
d�@|5�LzJ�	�R"c.���]U�9�<@u��X����[�.\�:׃v�z;�bD��@&�>�v�S/<!ۗ����[�҂Z'�0��_�"�6�Ð�XF,@2�TJ'xp���\�����"�nzg���`�P��v������>6�M���Ɓ���/e΃��qJ��􈑑�3BW�s8Gi�������|D��2Uw!�-�1�O����<ޥ<�)"��_ҁ88\S�/O�W��ѣZL�H=����g�Ύ�v�H�fa?5�T[�e�ɀzg~dgQ���׬8�oJHLf�粗A�u��:&�4 
,'�I�փz|�h�Z��|����:���3�v��b5N��*x��{ʏ���O+�fL��ǔ��o�9_�{Ge�s�0��N|��$���`��~+�f�W�0��BT�?W��B/ɍp�m��MM��V*�q��@G��$JjHxY#�?��u��ɉpV�5��� HXGŀY:;�0�ڡ��)�媂>ጳ�R9c�p���G���Ԭޟӄ�J���̌��r؋�HF111�2� �B���f���קh��s�ʼ<<Tp�"N�WLO��ٟW�p8[�Zۣ�n��^VV\�5.�����5N ����xHXu)@�M7d����k,�3 ����7��N���A=����wy�Ed���T!1�B�@�Ģ};#���j�0e�n (�z����xXY 2�t�o�G�2�?{&�m\�4���Q%��	"
}4
>��Ae{���tp�!�cI��ٳm3~�C��@��xR����]�;�����e�(V�"�4�O�l����/j���#��خD�T�'�k�Dpf��eTZ�OՌ���ݥ����@�P�kma����#�gE�醬sk.�G~Z��~���W��Bލ��	���rŤ��Z�+1��r4�u�=��4�ӟ%����\�A$�p	Liְ�;�}w	�8�On�s\�Mp%�aA���mU�@�wuNw�3B,�V%:����WX@RXS�p$�ܵ]|�>������7��:;�iF�-ѝ��qBB��	��|�Kxn���om�L��o����¯��._J_�iV�L�q�Vq�=��7.��.�B�VbRN "T��T�h�f2�t��	Eԧ��ZW9"h,��{J��(0N�����0bWI�ӞC�.�$�ԋ��*��Q��w��|�2|��1��n[�I�c�F��bZ��C�S�p9�<��\����I�Fb�##��v5aC�����l����"��������?+��|��ZU�;���k�[+)>)�
��%����?��pu�u�҄��ha�L>���F�r���KF|'�@%�D%5�$3�<o��X�h�����Sn���A������p��Щ�2\
1��;P��=R��s@���E)� {4wgg����h����������L�
�I�Z�.����(��<��Z��89���������~IS���6�(�yT�3�,~��3L&փc�&$�@1�;���۠�^�x�V]囻Lt\���0����w �Dק�z��B��M����.)��"�>�?5VH����ԑ�[^�ח�sձ�.��I�{��F�c[�h����w.BO���,I[G/�)�����q{ncк�VB��[�l�b�2V�To����(!��8�#�!_!k���
O���/â�8%1p��3�RD2��/�n�3�����bRyVc│�Gv@�f�xD�̹�HZ$"�1�!�9T�nڰaCSGR.U�Wo��^����?�I��y��b�0��Sj�&���o8!� �*nǭ���q#�� �W�1���Fz/���&D�\w�Kq��?��Ts���z��λ��iؓ`��$�q#9%�3}�-����X�߱;� W���L�]$����kP��G�z���:PX(��M�s�x�d�[P{@n�ש�á���l�;A�6��9(�Lݻ�W��TaK.<����E�i5�N���͎g���B�vac��w�]� ��x؅s&�)���\��NB�Q�n���{�x&qX�@V�,=����������$�5ڂ�%��5�8B���=n0\�i� ��44�T\�hm\��)�N�����O�MlQ�R��Vdu����	�/�=.Xx͌�Is��?p�*oHkjA�k���Q3�j3�Y������L,U���J2�A�wn�"u6�-ݥ#�OO:�MT��[�6�4���r�.K�绁����������ܯ�R���O�8�
�O��d�Z�;@�ۤ#-�������\L�mQ���8Ќ����/_.�V�����by[ >E����'��>���PF Q�Ym�#԰���{�4q��4*4��b��+���������;z�ӫ2A��Z������2Ϗo��@x)�~{�*f3, i ��	z�O��5�^���`+������kb�}��)ARZn1M�,�o�r��0���Ξ���y|||8�l%74 0�co�dw��&(���i��{7n�e�����-�����ຕ3��=5�N_H���]S�fe#��6g�Ί������\���_�$P����j}4�zR�.o��1;�Cz��,� �9�ɉS�k��G!�?}�t'=š�W�J�^��N�hF�j��AQ*���-�E�tO�m��r5�CͿ5�C�x��nF\'���#ߞBuզ�q��Ü�#�1�����~A��@l�u������!�¶�9]��W�<��i�|��M��'s#�ZD��{���t����y�U��1�4��Gihss3U�����7�9__A�a����j�2�L��p�ME�`2��wC���If�y��E�J/ �1������tΈ�Т���=q�`�6���\:���N5:s��T_����f,�^�G��188x�^��3��~KA4�g�[ �ַB�xp��p�$*���K�ꄼ�6��]�1��)�w�rp(Gb����7��¥�eq��a���h�A�=�f�z�u��R�7�̢L~�j�)gqɮ��,9�X�z������P�@�a��>�����~8�۞3�����Ɋ��K�U'ż�D_�Xxz�)�e;��GOx��]��l�i)�c+1���(��J��{$Wxu?^_��y���t��v8۞�߮1��/�}��5�����[����X�����*�vȫAQfc�ˁ_m�^�]i��|��qm�;�cU���2�e��&6�q]����ns����@8�8��_�j1Y�5��c���_p��kJw�B�/��(�Y����m�/}�}A���5ոSAkEd�Q½r��C{���3��,Sp�O�����%�]x϶z�8v��r�A|Ъs#?��;�ܢ��A'��0ޛo�?��bW�[Fs��FI�T�,A5D/�,س�D�jal)M�r=��ji�^�����t9��(P$�s��p+)��𨊁J�Y����}����.���qO���M��s�w@����[�������4�4Z�-}u�u�����6=v�u�D�k��ߩ����4�Mz�]Z.⁶5N�3���YX��6���r ���->)G/����&�-S�gE�����^mWp�Ԍ�\�&{���!��FX)s��p�e�����z��&�^�̹�nӈ��Ϡ6f�tv�;��}lMGȔ%AE�q� aO�+��\]^Q�_�Ը��g�(~O[zow���sLs�Y�����r�K������4B�E�	��ȇ��A}}�--v4>[{��h�6�_W�%�6sDO���І/҂"�d4���((n� �L������'�k:"/�q�����H�8�}���	��؈%i�;O����h4������߾��_0{�\��+*j���*�T���0u���lf���;�����R�\���Tuhί�'�>��>�
O=���������ر�3���������u���?j�r[�`�|z��X��L���^@�9�2�w�ᕪ��E�5I&��i<DX:�ܻg��S+667c�[�{~լh���>�ۼ�U�?�.�=N�k\s��(���I5��|S�vn�����V;��*����1�ڗ���8�y�J���7���^9���O���|�Q��V�t�˾*�T �r��cu"%zžt����#.��u�I��ǳ�f�1����Q��^�5��j ������s���fFF��Kψ�Yh�m|:��.������VE�����o��Yv�l�?<���M� ��ǝ=;�D���6<z�䬼����oW�(Kn�k��)��:�0.�:9��8 �b,!�0�(��.
H�^�d�B�g<ޗmjA��� w�q�1�����eO?�~�va�F�m��͟#7{��@��ƙ��G�q���7Wnd�_r4�&,#�W��h��8_u�b`as�K��>i����3��ܟB��=��R��&��|/w�Ϥ������Ig��5-���"Z_ed ,*j ,~}���4���vۯ����}=��ā�yR���`~lsNϟ	/�ˆ�H�x8�a��G��6�*�o?
�� ��q��#@w�F�c"�������Oi;Z��rf���ڗ�|eD��㊃J/`��JD�̀���Z9��V���c �x��q�{�vһ�L��O�ܞ�N�܅�_��z��[���!侲�� h�J(#�\������ં8���}�� �F� �����/s����r��LS>�ǣ��酬6�� \1p��+x��U��A���v��͊��2���g<��C�E�)w��u�cGj�x��=�8q��y{�՘�8[[[-+K{v�?��V��I;��WrB]I�x~���.o��� 	�f1g1.W�mZTMm9�� *��A�W��G1���q���r���;�M�`�N��9�C�n�)3=�ԴC=���!��:w�A������1����]��!�t6⡴^�k}����0v~��;a(ZNc0���Kҙ���Ofi.�ky�j
�Z�}is�ʘ��͊���.�|���e���p�O<Q�������Ui�
�:���>Fl�N�dv�D��#'���Y}B�Y����Ļ;y�tR��oI��j�^�ۍ)�@5�]�T[Sw�O>�٤�!���?�Lln6�R��,�_5��H'''s�YĿ�W���V'��b���n��)c�mq<��O�����!-�ǌ�ה������
�D���:3�t���z��mn���Q�~#j�'��b�yK���L���
�����sz�lc�e3��E�Q�w�e����e����g�ƍxnh�+~!>~�U���P�b�]�����hy��P7�/�bG��|̂{���C�$��9[j[�߸��_����E��s%�N&��b��h/�ъ��y3&2�L���C��>����&�~R�����v��Zj��x����Ö@�r��v,����fE��/m�p�zs�{�ܱ��Um�$9=�/��."�|���TXc�����}�Wq����y۩G��@����-���/;�xAj�M�j��T��N�6�!c��|tH�a��C�!���,�U��*=���!Aתj�'����m��M��q��"pZ��a�{�j�̃�z�ϝ �����TӁ؊����Z��(���w]�,����/��ܶ >S�������j�� ���=�S|�����..h�fp?ah	�o�,�K0nb�/�`�x�m�(��EV�3�bEӌ��X,�se�D .��%wd�q��k�׺��R�:�/��$T���vA�����CwZ3n��t��/=wM�9� ��鶛+���2z�L5��)G	�\���5��O�ʫ��U9f�3y �3�:�o%���~�x8*k)E�X=�[\����8���{����]�z�K�-�=��\N� -xrz+r+����}=hM���Y��4���.1�8��\��$�5_ͨy���M��ŝ���#���x��	��Q|�و��΂�Z���P~�~�N#|φJ�2��[YY)oق;K?X��`T%���x2����r���P	���p?PXZR�������������p��V*�:����?ȑ�3���F̍�u&`Ѹ��^�H.�nqb��g0���hX�&����?$�~i���(������ᤐ1uƁb��"���H�ۗ6P�
�?hq,�y�g�	�(\^�0��żlѳxl����b 2���s&'< �n�,n�S���3P���z���a��l��2K}(�_�V������Y3�C�-����q�kfB��	�i[l�w��5�ʓ����K_���=�vχR�\�]W�����e��&��������LP)�@��W��BM �8WO�F=8�Er �@u�O��/6yTՆ|��1���P����$��HlUՐo��o��o� ��+���sm%���^�(��fi��#�J�<�j��>E}��V��
4�] r񢟪As�{w _�m�	S���g�g)@rW@�9� �.��1���>���;:N0W-F�� �݊D�%@P|/����������O@�.��z6+�l�V�!�Y2�}�_�"b�~��0�II*qoX���T�%�������[��k�*��,]�"�Z_> vlºc:�b�d(KP�j~A��!�y�$�܏'囚f��O{�ZCN3��Xy��ޕ�W�[l쳺7[�w�.JFB��^�a��N���Z���42���%��iR��B��_4���.T�uD��`Zf�k�鷜M�r=�<[c��ڶ�g6��Y�!��l9U3���LL����=����Q}d�N������x������S��x �b*b���Ο��|;��6JM��p]�4�a'H���Wݚ%"G#���eD<��W�XS eN���A�:�����}�	�� ���.70)��P{%9��x6u��#��:@r��|��ضC����A�D�a�]�Em����/��M�	�`� i��Χ�<��/�H�#����)�����MK�l�8
>��;O*�^��hD�����e\���D�i���#T�抽�e������Cq����Eۂ�$^����+Y�����S<@~ߦ�
$A�Y�%�(��jm��i�B	��d��:�T�2��D�S���%�Pl	�����s��,q�Ѡ"�1N��P(/}5?6rk�Z�G��'�9�ف�WP�("��&E��l��)��gl��>��##O'~
�� .g�?�d�G�Qx���)wۄMe�3�M�H�$�/��O9�$ǉ3�1��+O�TfZg���~훱��N�G�JD_q����΀���{�K��_�>�m�~�q A ˋ.�Qi��7hl�n(K�����f~q�E�Ts�:��|��sU��j9#���{�R�����J�u�bn�΍%υy|���8���޴��3>�����57\���S"�2�z�^zb0�������&e��Ε��4��������j@��W�p<�ǌo�mT�k\�
f3��ջ���MoLq�=�[���ij{
�HNR���2�����<�@��i�G	ml[Z-���ك=�x�r�?8����ZN�f5dmՇLNe;=Tax\��5�Ew'��[DD�!p�_�h#���?m�p���SG����D�%�I���o���hS�"�$���/��8ٳlu�� �� ����Ӑ�S�X��A���	>YΖ��L�ZQ<ػTY\�l�=sx���g����SU_z9�����>�jE���9���������?0��3���E�E���@J2�"h&������.ǀL�� �p[�S�o��1�1r��P�@Q�+=�:�[����E)t0�$[)0J��|���(����m�J�?���T8�np����������g�������ˬ��|Q��~ b;�\�ʠS��K��J} 6-�9�g�>US���^%h���Ӫ���s���na<�Թ��YEE����*�7v�]���;�6)�}����f8 z���]9��_�R�f�*!���l�]��W�6mmE��y�6�6�%��֕ ���
DI�ۋ﬈T?�������]�j�{����Y�� _�����>e����4H��&I��h��'�{C������\��}M��Of���<�*��1 ,sO��5qA��PH�r��)��s{��3�$5I&aω�rqFZ_���jN �]lmUܞ�sZQ�	��F�S�rX9�i�2��b3E6�@^�b,V'r͵?,cڜ_���M"c��㪭��Y�� Q��P�8�c��i�w�Q»!/�rxm�#/ԟK�<�`���������)���Q�h����7��^����,]�z�^�֫:\�x�>� ��D�̥n�YXްaË�������땨�|ųjk�3c�� �O�/�g�/?�T���pvOc���sQ�s�(p��V����{������,�<ŊT�}�����ݬ��}l�j����| 6�Tm�Q"�v+w��|���ZJ��ʓ������o�n������!i�Q��?|�z��GskA�WN}7�t>�Ε)r XN_���P�A� 8�ԽvT�|/��?�+�zl
�� Aa��x]�����5�`3�6�Uye� �����c�`�ZГ�2������ӧ$�ief��_ �8�^r���x����K�P��j�t�����<�~��uy��e/��9,�h*�IRR��t�9X*_�b����C[���BR�ρ� M��hP���f�y�v�^��Z����=Z��;�Iq3�hP*)�KQZGv��yj,^$k����L����Txӫ���w��	<C҇���ƍxmO�۴Ӹ�+IW� *���0���-����~7�ce�TB��]x�ů���G�yɧ��}�р��6N�M�)ՠ'.� _ײ��%��/�UV����5-�XVԪ"~��jn6/ku�X��T�PR���2$ݾ��ݚ���{�>}�I�����Q�۪ؤ��B5Ȫ�3o����N�0��0�l�6�@�a��!�Zi�w:^��?�ߑ*����?��c���j d�K��f��M�N_��[}�ˏ�O�����R&�Gn�Zq�Y��`n!� �������� �� ��	���c�O0�:)��S��ۙ��)q(b)��|�Ry�gf��#�DL3��5���,�/V���I�v��X��G��A!�zp#�V�?!��=����l��O������k�}^�k�r���a�g�0�Mw����8�7�'�Ó �����6�!Q���o�$��c6��3A~��t��f�C�; ĝΩ�ܝ����
�.Ew̋�ƭ�c0Q�No��A�سŋ*�U?z��X��2�w��D�yaP�V �'&%�	q=�4g�+�N������d��D�E�B��e_� W]�`��Z⪛��T*��� L���b�ʥѫ-e��]w@�@��i�:t(&���Ֆ��AAH�"�sOh��G�=� "_[Gg_,�j�.�IT`x)������05"A����Gb�ӛ��hҮ�lj	��$�ާ�I�=��s���D�Z�eJ�	ٯ<�X��窇��|O��oe��<��&�Sg�����n�F1��@�u�<S[�l�JlcO|cOǷo��ڿ��õ�zk���+��|��潐jڱQ`k$@|,	����&S�e�&��!vA����j�Ԅ�W���#����6����	�/W�Z���v���Kћq�e�c�B$�rZ��(�[��x&00r�""�����kkkC!�k.���`�وӔ0�ƃ��o��ۇu��62�P���P��GNk���t���9�4�T]� K���o�e��w�5s=Un8*`x����]p���������W�q;�d8@�"OMM�c���E@����j�"�$�c!�f/��Ó������n��˗���E�3)Zn1Ne*��==��V��%܉�0(ԋ))r��pꔙ���/��4��j��!}���8�d~�έhF�)�,u?��B�����j��j������&�6�9}0w��1�R� ͘��)�
D��N��;�%"��	$������dS��?֩�@�@Qn2�,�Y��36g����z��́��L�5+���Bb�MCmjz��
o�1(��En�J ����?���	�ʂ��m�l�)σ?���s
�Y�1���x�ef��Y�U���������׌h�W�X�����V7�g��R��d{�ԁ-�Q��qF�%-z�΃�D(��VTT!����g)�>&�!� �:+	��#�`m8���|
VΥVk��ws�ۤ����h�����ZL���9/��,���sx��v,Uq�=�C�v����I �H��m���T.����5�F�y��z�<W������I�-&�ꘉ:~�{V���;qğ�sj����џ���Q�rl�Ǡ�>H������@����1��ڜ��ǯ��m>Gbu�U*1+w��_�{��و)Z�}�����u�R"9���=��69�;E'Y�.�K3�O�>��I���?@��VU�W26B���5����z[(��f��cc��k*�����39<|<�ء���^=�z<R�v}k�WA���7}j"��p0��;��-�:� 
�pLm�ȊV��[�d
�����c��l�Pao�H�e;��)ۃުqV>l��k����NՁ�_:��ZXV����C��w��rW�9;���C�� K䫼��yN���z
�M�iM�?�^F/Tk�Q^�x��=�5��^Av��\������%�~y�0�^4L�y�����75�q&�/z	���Q	E�4��A�û��و//Sx�[Q�3�K��5%��>��qͮ,����8��c�ɛ��!7W����h�O��ɴZj-��,�g�G�^5ejG̰�2��y)3e��q��y���Z��8��Zv��1u��Q��<�vH���>)�k��Z@]۷i�/���
���0���T�_� ��(}^�H�ׂ��:k�<����~*������Z�iYP��KnV�<s��jN���\��+xeq�`�BX�e�gu�����7W����A��R`'�E�7�������V�lW������ì�L�]8�{�_ ݁�>�~�ח�S��<3<����
�Y5Ŋ�S��[�.���E�!�'�ovt��s�]_"��=��G~m��~@��)��ޙ@��K�ǃY��-.@Uq����T7�6����Iҍ��s[���O�no@�V��#�����]~/_V��f�6+�Ֆド����?�v�g��ؗ�0��f�gWcP
��,�Z����B�9��V��2n_��`��
ϝ��{Yk,����a�3���a�`������r壦��u{�U5���#��aabU����,��Dq���,Ӆ���0�8Q��:P�{e1��غ\I��%g
���/�S��of���cO%9�NrW���v�{���_x��2*�$g~{�����QM^_�/�`����H��R���J!@UQQQQ�JQQ��!j+
E*TP��+�yH�H-j�h�!�m������������w׺w}�X�&g�ó�g������N�*�$y����7�Qsm7�bfi���w�?CR�/`m��L&/O��.�.>X����R���vIҝ]N�mk�izSސ��J��-���«Ι}H�v�m��C�ba�)6�|:�,&�ԷG�5���Ϧz�y��U�J��)�6�|��*QG��km ꀅaCe���*]�X�h��5��X�i�o�\Q�l6�V������~�hƤ|�%��E�rY����-��g��Ws�[�}m{�W�eCp	J�eL��o5�"��%7��_s2��6KA��ϝ��%:�i�y�b)�Z{=�j�cGk�/K~���.{%)`>��H��.ٰ�8JՄ�.��/i�us�_{޼y�ʟ;yb�K�٥3f�4���(���"�?��tX��*�e�p��A�Q���>0���C�7��H����ԇ����M/:�\����yr �|�$�	hR�@�L�M��d��:�P����MV�F9�!�#��AƆ���(�<�M�`Gxi���+򍐷0�8� o,,���7n��=/��S��ϟ_xcx~dV�jI%�@䓬�R��&��A][`�`����>�9�-��S��M#�>Tl�h���m�a��? �ݴ���z�{�e�@%2I�M�펶�>���@7؉���1x�n/9���� '���o���mk��`llLs��ӯ�}�G�]��	����%Z�Kc���K;E�%�; |�E~�����{j���to��l��f��SK�|�t���Ktzq�����B�+�:�<Mt�c������{ףΆT .Dz���;�!!%���g\@ۅ��C�2Z� �@g�xa����������F��l�b��U���b����6��9���P�B��\v�*��RȤ����I�����-�[Г�K0ua�N�	r�m��g���/�_���B8������P�㡼Tĸ��-�D�1�wǷڍ�7,G�ƫǎ��H%��Y�c+�S�(u5ꕲ���a;�#��rU/��aT�&�턼�Ps�٥�Č�۱�7�����d�8p�Ӛ��>���p/��Y�*�����;#~<ඕ�b�)u�e�p{w�7W�6V�
�j��u=xt��I6c�_����'�<��>5����~��W�u�
���CT�6�:m���(�j����})}�g��� �i^���Z*/Z�YK���#��%��o.#�����pD�Y[�GI�T�����%f��+̃.z� ��*Lj^���n"GRϕ'��L#J��,t�F�Z���f_�L�'�����gP�::.M�Ah7����Ú������Z)�OF�l;��ӣ���*�����fHV����~����]!��{#֒���N<�گ����|',"�J;M�Ɖ�~ŭe9�%��(�[���B_��嶔_1?1������6������¼���F;��M��Y��>>�h"��Z����U�0mM>�Z'�cU]���z��hp �~��#������\�q#��
������NN�V���1+2��-����6���ۖ�I�� �2R&9s;�4�\׀�o�����]�s*/E���,�v�<�&� �����a88!�6*�/��L>�6 �/�ҷ#�z����j#xF��j�����qS�B����:_rt:��=qx�-ϛ��>'B�P�&th�-D��k?OŜ;��P{A�]=v��C@e��A�G�Uȫ"�i�����(���6��g��P�B`�/��Tn���y��5��ݲ����Ɩ��[$��C�F�k��2�8#�Y�O*}�C�����Kj�E���B�}T�I�C�P�Z)θ���J�F�=���r�Br,�i+r}Uϸm�y��I�����<�v���9f�؍�9@%���bU37 mT��7��+�&�����X�+W��]-^�+���7���f.�h	����Dii���@)�;�t��q#n���>���KH�E��X�`V<os�����Ď���p��ze�)��Jaǟ�u$Y��{�n����6A�<�c ���ϖ�a���/�ʆ��H��ub7%uɕ�;SX�^����s�>�'g5/M�����"���m�je�7��𳀉��Zό��J����@h[O�\t֤�BC^O���sj*x�ä��ȯ��"fr����tȫ��bOǆ*-�!ƫۤ��Oоz��#_��HN����1��� Z���@��*�|(���}7�g�����%����#��\�BQ�f��m%K�p�@�"u�����&W'V-8�_�#�_{��gA�n����`�����.�q�� �0���,�߇S�[�<��C
i�/Y5&���:��K8`( ��տ��[��x}@W��l���¡����˽6�3��wGj��/1^��Zi�L���y�=��x4�=w��{~�=r��K�g��[������з�7^��ٜӉ=	Y��uŊ�׿?52V��hj[pp̷�Ϭ�$����5�W��@鲄M_��.��w;�X�9�{>��j��@7�s M��M -�����j��Z�l�:��6�!��K}�����У]�.�D���<<<�v�٠���ܒ��4�ʫ�o�
v<X�+
�Dgo�~<�{�����7_o��r�H}Yf��݉�Ve��Il愗7����
�Ƌ7�C0�;�4U�%{�S
���.��T������E�È�\/i�c��2���;)R@-x�Y�9v����N��=�.�g2`��V�ߪsPC@�A���5�ҷ��ŭ`/ד%���5��1Ͳrz��HqPŞ<��|>�?��O�b�|e��8#�L�ߦ��_���o��!(#u��#G������Ė���B\F1rk�,�����d�5�] �<R	��Ú��eD�R�*F�G�斧�����O�KԜ������aM��I�h���%�|/��Iw��t��_<i��2F�������Ww�}̖SK��De��z_�����XX�f��oL֮�/���F�;�aD��y$SJ�N���v~}�;���f�h�e��tI�d鄰An���*_����v	��ߕ_f��̛{���[!����4��P,���i�8���ޡ�r��e�&�w�}����G:�5\�z�N̍��}�'i{9A��_~#(L���O�X\���mv�(�a�A��y*���ſ.3�U���;]|��8̹�Y����"�մ.�0.����.`�S���u���[����zB_��Z�^�s���d��$�����[����$��rb��P���pM8����ymA��QҺ_��2ys��=l��囼(�-//��!�w��*ݰ��͎��>�
#V��_����K�Q�~ӜL2�Oq���_�v|���E�VC=Vy~^�i�(-��b���(���B��M��_\?�.�n}wh���e~�A�r��Eׅ��q����s��TL�+"`�	���3}�}�e����eSbl��b����&:��[|��a_a�cS��W{�ND{j\�Ζ��
�ߓK�Z�}n��v7�� p �Z^SW�h��NxF��ih�jg��`�L�����w�,��九]]�ys�{$u�� �;D��=���)�|�����b���nm�e�)pWM��H[��8X�b^r�Z�r������p���"  �m��!�2���D��q�lEߎ�>���4�R��0˸{;�G��c�� |��u�B���yÜ��0��/�mg�� ��*�A�G���M`w���N�����oG*�B ?%�?�ΰ��/\�?����_�����>
���/��D'�e��`��e)!C���HV>���g`<�%/�!���g��+m���]���̡+��㑒�9�'lRk�@d5��߻�X99�48L7���m��MM\�"�g^۶\��4:+b T�5&O���M`���킙��{����h+�A\fT�r�A[�6�)J]a�əO��M����;�؝U�Q�`��,}��1���o����Y][��a�n�U����d��k�&����B�z8X ����5�٠�%��K���v�`���OM:rs�����&�Q��L����8�M�dmX�V�2{p����?��Z��-�g��g+�$���rݙQ�_,$v����(�ͱ��Z��v�1�Y�0�+Vf<1TtEr��c�R-�+'��������p�w�N��a���UǦ��8��7���N�� �`_!<Fx8�RM��z�����cJۇ���@P�⏮0��	I�C�<�4&�Fs��9)���6q|�E9�T�7�MO�qҰ ��RFcMnd�z1��;�N)�ώ��&^���j轣n��� �P�:4�VXN~�� �=wTcΓ=�������?�"W�[��o��Yl���:�����l[(�
v
Ѳ�ҝ�y�A�n���wr�(�����I�;�	�;�,�s^OMP!�ّq�X����_�l�4��("��YC���cK�%q2�%���e19b�M� �[�M�qu��D*z��$�-�:��wK$�b�������%U��D�a��ی'�Tg��k��_c��*�x/vA�,�A����N�zXKS�E�W#��R׾[r�Y� I&��銣n�s��P����@��7`�!	#�`y�?���eS��3ٽhR�e�%�M�	)�� �ao�&�Xt����A��-d�~�E�����C�
<�ݬ�u5�,C<�D܁`?1=v��]�077iG�a�kGS��������`��zBS��V��jM�Y�v�7T�-�����_�\��B U��5G\R^�oE��?��0��9v�oL�ж��p�����g�3�C�G��ۃʷ%ǯ�KN7�\)6K:�2X�������s@E��/>:�7��_Wm3|y�T�b��6ggL�
+&@�=#���>:v�u'�M��3����'�
RY��d<�|\n�Q}o�2�J� ��yG1�U��-}"��~U끍�����E� ���2j`Y��#��8"�ڰY��i����U@$ ����;��Ի�J@&� \��Y�7���=�*��)�=�*��]���:b�d�\��oq��-�bs�/�X��eb?ў�=؛;oj�@���7�ᛟ3�\��M�M5,�r�Ż���%I�E�[��^��"F�;p��ܩ��giF���=��\FP��nC�:��3�9�:J�}�G��a��x�:�9!��@8�C���l��KH7ع,��ԐZW��L���n?z�b%
�v���e7���u����o�EA��]��c�oqvxߖ�����2XT>�f<X�������f��#v��3`��]�@o�ZnSΖtО)��ҹb.��DS2(���w�TF�5��T�I�\"I��S8x:U�e&'7^*���d�ذ�c��V�� A��])0}��q�ug n�U#�bt�����YQ��v��za\xzA��	��a����>����Ď�z�X���\��,C�[gP%ΐ���
-�"���.�cE��������'�+�?C�����s�ԽZ^A�m�&̡8�m�C�[	@̶�C:����7aX�4�Lu�^�����F�\�jT��/��{�ʧ08�>*�Ԁ���le#}n͹"�[�Ű�;2!`U��]r�4�4^�k�t�)�y�~������4;;Z��d�g(X�{���<o�Ob���+�#��ZS�Ȟ?������Ƕ]�(�, �/1�����ȜSsKb�N���$��u�'� |�S�+,�2*� �猤�3�:��)�Fꈪ��j\��U`��@��Ϝ�1�I`�(/�{O�v���E\�����Ȍ��Gm=�u*�$`�ڱ�W���	�D�8d!:�v��<(��B��p@epC��g��Γ�R������&�!�; �-QA�H�Y\֙ч)��	�����Hs vŲ{��P�O��G��� oӊZ3A�T	;�\�Pײ�S���N�������J��%� �&��p�B��ݻ�K���
�� h���	T�FP�5���e9r��	�+7×�ؤ�3 ;��H�&�d��*i��Ԯ&��2�\�D�'E���
��K]SGv	��_R�'M�3rĎ;	��q���� M��Hp`j.�K�8`x%?ba"�w��[v�'��LX��b!8h\�*G�frf�߶:��7�ĎG�U��F��c�����y��7@�%}=�(Fh?0�]��wM���`z�{�WT���z{�������+��N�ķ�TУ_�����ˋ�
�
ր2X�,��H5�B�r��U���XP���h��u��P�k��kS3�)CyT2�D@��Ď��؃�`o��v��M(�
*��NS�>�j�1�����=�m}q)%;��W�;�e�(�<�U�t�N���<W�:�����e��{1]��.:̿٧R��;^���o�>�5΂��ps-� �E�t$�1�Q�Eܸ�#ª����PO���׻���3��0f�:`��V9�Z���\��p��7�Je-,"bB�N�-�4�*	������v.g+VK�*�T7�5<r@�c	bhoP���nDx�a0hI5��(9sVh��4��� c�n���0�Ŋ6���	�4���ٽ��X�]@==��$1{RL�ƛ�5���!�a\�dM-���d��4�
	�/'h�o��hH���.�C�WL#F>�"	 A���Q���y��YU�a�k�N1��`LP���q`C�W��}�Һ��W��D\�6���@��nѹ�%=�>�*��*��+fp۽]V��r��J%k�|���@���b�=��A(�R�^�Y����d#zK!�Ĩ�g��oG�_A3QE��� p�x�d&�M�턄��0��j&��BST�#���I .>�����X��n���9�ږsSU�7��,�G��k$��k@^�� 5>ħ�Do¢uRc�����-_z���BG$t�����'n�2Y�V0J��4��J���f<����>�;��+��d�E5������K&^*ۧi��v`i��|C�^\��ȁ	Tcѿ?���J	��B�#����s�R�R�&��Q�/���Y��a+%���o���K�9�#Ek/wj���:k�C툸6�t=�((�Ԋ|�-�!��C�r����1�o�=$'u\���V3������U�Q��_��g��Ða��c^ ���ư�6 ��<�߶e�6;fm�;�ߪJ#��Ҁ�*�wnҟ[q�W����i�{!�'oJl�rF�hMM��� �E�)���b,k��;e5�o��շ��34�n�bq�i���U��P�jз3(fܿ�	UN����
��
�D�4��\�.޲Z1%�K�%a��+��_��5^�W���+8��v�K�O�&6��`��y)��}����h1�=`+$;Z�s����0Ki���ݲj�Ё5C����I�v������|6��g��f����(�C7`�ITl$�!;�!� $:�t���K�~����`�.�������e�i�P݇iY���^/ˈ�-��zNe����Ņ���;�H��߲ҽ����Ô(�ɣf�ф�
.q�gE����B��%�5� âw-�
��m�<���޿����K��T9cR1�8������`�'����v.{Cj�����B��V��T;��.%j�[�ʌ'{h3��(�擼��C��P��6!k^�#���h���XGPY�lμ?����
��Gf���+4~1��V!Tou㸀����������3}��~.,�P~���$ؗ ��N���i�����CZo�FM�b�B���9��9M���cE �ǚN�5k���Ո�VǢIf�J_\�*w�o��Do��������޻d-�/HA๶x��]/�	�4�D�J�4��p�_	��xql�dS�Ѐ�x,�|�x40u�=_;�[�!�J6�v�UXm�o���v�eX1�r�8�u��S�G0P�&�T� o.�B�"��m9 q���.^b<	��|�L�~z��M����c�s��c�:��M���G��͇q�4��=Bw+�̯p b�WJh*B�^�e� �m+���k�kK֑�h5Hi{�5��v�a7��L�Xe�2"w^ M�!�p�$�<ܕSF��j;�^��d���Ī.��P��I�T�s�˓/�Sd����f���駲{e��#�g`�@"��Y[�Kҿ(
���X��?tO�C3jQ�n�8L�Y�P3 ��&�x8�T{�tT�xJ��ى�� X���%��1Iݦ/�b��<]��X����u�vL���Y�/��Іpď"�J�',.��������aM>dߢ��u���LeH̺8�1\��u�6�Q��,�"��H3RZ V��)�����n�!���b��^�!-R��uHq���GПf� zHF���uw��>��,NX4��=$�E񲳳�e�w������v�s�.��$eR�|F&�璈�3��Qw��5�q[��%m>�K��+��؅��Z�f�1���"5��1 |���$~n���H��D�d��b��WÔ8 � ���͑L���̚3����@�#���w�#=N�l<�����U�"�]!"�=Wz���B�]v�D���9~��/@�uva�A��� ��b!��}Q��|�
z2 �6��"�}l�v����\! �C;w��ͼ��Ǔ�^ w�Wq,
�����N�}���C ~xOtu�d�p;�-�@q�"(G���{��)�. �>��NS�8�%��<��'�"�1����iҢ����8 d��H$dǇ#L��<XI�_@�Ao�����bpz�Vg��aX#���L����ؔ�t�o������@��I��-W�O<=H�#�Y*9��# EY�g�@`�w���*��&�'����HnN ��LeV��-d��A��}�(U�x.�Fxeu�$�i���?2��\�%�L�#��L7
���5�݃]��D&��&�]��~b�L��Y�DX�{��Ws�a%�����!�F)f�&�5M�N<c�M��.���S/�����A�b�2�Y��9����\S�����^��j}�0g�-	�
T��K���&^�0���`�zz��i�X;82\B,��o��D���(95�g�MO����V�;��'�v�:9+M��� i�&8�4eI[=d���S�����l9��ڨ����'�͢'[������L=ym8�Fy���P�A���w5��G&�"L׆������1b�p��e���x�8�T��)����cDKhK��(�Vw5bA��<��Ԧ�A��3ؤ���C ��8���p 9�]s��\l�������6�h?�����_Ǐ�	I	{N.R���}�5���*��b��r�K��� |:�m�:����{�@E�A{�� ����z���g��~R/��0��EΞ7��D�H��ש|	��-Q��\�/����2��/6w��MPH�E1h[Jl�m�N��慸ސn��e99�k�\��c�a.y��RQ^Ԋn�s'�2*�U��=�b3(�$Gs��' t�v紾���P
�������Q�6��q��t~r7%z�A���.Î��&z���	�Q<��y�p9�+W���|���!.^67���>��M�l,�l��
���s��
A̟�b�t���$��R��=9s�Nl�e���]Տ�/�����Y��#~y����!l!�c���D'�힂-��&ǈ��xځ�,Μ������(Ѥ8���v:�n�n�	�y�ZϤ�1~Ľ%���J3�h��׷�d<�����z��n}yu��M"l���N�&
�v?����1�1��R!�OM:f_-/7ǃ��������<�D�P��zP8lyA�+�X�
"��?�?��hђ�W|!�7�Zkm�^,�m.�����&�3�]FS(o�P��,�$z��ǀ�0��^҇6,.���0}��z�����n�kvi��]�c�] #D�Lρ�^|���d���,���K�
g��� ��AMtk�}4%	�O�"��;$g��ߐP�Ҁ��5�^��we��
�eX�/n��Ǆ�b�ۢc��[U�g3}`L�Qތ8�[��S�IDk)V3�('f�Զ��0�9�q��� 辀�@�ȁ�B���5�?���N5�1yi���/��b�0`f�I�wYgڡ���f�\�0$mTC�qX+=��V5u�ЍW�X���.~p����i��}�Y�_A��L�+=��4 2����[��.�?E�� �N�қ4s������&^[k�
���N��qA��<d&/�9+ɀ��{πݻ��w�25�Ϩ
�8��}��<��P���|*�����zjN��Է���7�K�Q	�l:�E����ǹWz��FEE!
|5����T���\w�!��=�� ���՘p��s����I��B�i���g�]��)���򰕮��P���H���$�n�˝y�i�� � '�0�ۜ�I�y���`�O�@��̡*�}�#&�%yO�$���h
C�������0K.6�+��r܎�(�`&9+p�d3��	�l-'A���%�<���TW�D�L�v��Ut��C7|f�ri2?R���	mZQwD��qU��)������J����r$��Q9�aAM�=�:¬�i�#��5\�JI��U�Gľ���8NL;��;�-����E��a3�Rp��Q��h��Wv�Aލ�!.�K��[P�N�J�9ޖ�[�ď�S�)���|KW^��}��Mqj�[���:,�V���J�6�%/rǀf@�S��	P
��:$h+4	i�D���׻�w׽V��}sx[�� ö=�8?��+�s��m:̈GK#�d��!����a�wx�`7ʑy�:)�,mג/���cc�eZ�kD�@�����,h(��w�����5dl�'�p�]n��Ȱ�d��\��p�]z��PT�:%(�7:��8�ޗ%�c�C�s��c%� R߹��o�J�A,#*�7@E�� ����_P�n�{���0=%:v�-77R�������=���!s��úǄY�|�й9@ɶ����� Uc��}+(PP�|�RW��iV�E�<��F��y���U��{b� ��|�+Z(S�?-��7�yÐ��~�{7��{�b�893����!Y/���J��q>��}�3ai*ƾlnսj��|Ȉ~N�3�cj֬Y��5|��tYv\�nUdg�U�}ﺽ{��!�/yZ��s�����;��a�����#̦�u�<<"��M�8-!/lT�m�gT��{~{�ഴ�qRM�����I5W#��Z�M�♧�XI��]��=n?�3���
�����U�.;��l�)��2�PE�U�߇��{�ݎCn��g-ѳ��J#x����WD��)-��rY��������d�r*�'d�2�蟊�J��?�J֣�1�;(��TZws��g�2�GP�UV߿�QT6z�yഗS֯P�X������oL�>z�����M��2.���<�~��r��'>��3��W1A��%�k��5K>��YO9�/n��H�|s��ǋ�4�G�]�-�]R��ݝ���� �U�C 0�����'{�322�PRy�q�-qYDeII���)_��v����h�t�ewV��#�<|�9KT��t���a-}��Gq�]A-����m������4�	?M�i���6{~���o#�I�)Q�Kb�vK3����5�j}K>���9555n�#�-�a�ß�KKT������}w}4:����*gi�R�����mK�l�74N�]Z�J��?��?�WMZ� �(�����P���?F�_���mnܷ����i�O~��ӄ�&�4�	?M�i�O�wZ	�H|����Z']2���O��ѧG�}z����(����%ǻ �/��ӣO�>=���ӣ�ۏT���\��>��q��Y�y�PK   �rZ�GDU7� �� /   images/d628d844-ce42-4e82-be63-f5fdfa438334.png�wTTٷ.Z6ݢ�@w+���6�d$g[D$�䌒s��
[��,Qr�PD%I���"�Ud(
��Cy��w����1�p��[ٵ֚�ߜ+P��T�~��+�����1q����u�,��oT���g�����{��%���Ώ�����3-6������k8Y�#��Z �H$������gn'W�D��5�O����5���?�9t	��T�;N���h?ڏ���h?ڏ���h?ڏ���h?���-`�9����t졚֏���h?ڏ���h?ڏ���h?ڏ���h�W�����w�>�d��c̯��nq�������\<W�^�)�����WvK��[���<���N��s����vK`_���jv�z�n�����[�o��p3�=E;G�oZU�y#3�{��4�.�����o$��0�5"���x���ȏ���h?ڏ���h?���Vh^���a=)n�$�pX޿���g�\�+S�(�6��](Ӏ	�N㱒�w�'ӪJ�����K!�:Z#�|��fXN�Ĳ�_���F�cv�n�|�؝v��T��m�"���2��/�r�f
y���f��XH����S�V����z��y!�R/󘭮3���g��o �3����Z]fk�>�)IN���;���n>����9�}M_iX�X
$��D���������+��\����4�ͩ<Ƨ4Ƨ���)?�Բ��W�`T�SY�V��o�j���$������eObՕ\���Ն'�k���_��_*K���5�\��ubK$��G�0 ƓT�g �\���	��i5O<�yfMQ
%��ޛȻ�T�����ښDq���F�{L�ڈVav��>Z�f���Ԑ���dC��^��?���~����~Z=Ͽ��%.�
�d��m�%����_�)��$��e�9��LM��#����s>s����4Ҩ�S�n{��)���i)���;�z�ֈv(�]sh!:�v��|7����e?�o��O{�'�T$!Ћ3b�V@^n;^Z��K^~_jҤO{j�/kM���u�<+F�K��)��{yY�T�������^0��,Sy�/x1j�N`!�X��6'C�c!sB�]����E=	��CMf��]:퍹����jؤ�gq��c<�����Q��.V�Ϣ�e�C�J�TʌquoA���Gs�������3�9-C�퍽.��>�ٞc�}���E�'���q���~gJ��^,�)G�M�O=&KyA,�$k5�呕�������.���5�9�Ӹ�?��6 �jf�����5��� ���˔��l�2[���	x���r����!-y�79'�f(K��Ȉ�cl�� ������]�R�?�g��EW�󝲯�l�]��B���(�	Q[�%h�yM^X����/{�kF���Xy�ZӤ|*p�W=~�
k����N��s�?*�K�.?.�KGi���>4��w��r
�C�'�8ܖb��W���Ȝ"iIS������)�3���/�c�^ֿ�����?�;�,XF
��ߋ�T�:e�b2`ȴÏE�n�m����.	��Y�Cj-S}�22���k��ͬp��@8A�(^Z߼-�H����$u�l�rg�a��,�:2#�'6���ϭ|��j��^�>��=�G�O)�*Yf��mڎ���FT���)CM��4Ly�'���>G�=:Iqc�0N����M��9{��I~Sf'�߅�=�WV=�,�9��Bed�H��Hbל���KN�%{_/����bo<��K�X��0n��U�����}��8f��
h{�춡+1#�f����Q��!Y� �!�~9/{
V2�����qK
n���X8<�#(c�!(O��m�G
� x<׎���������W���Q��T;4�����3���~6HB���ۄo�.��BF8�l�0��ܹ��G�d]y,��Q�Gx��8�oVSR(>'��q}�%�"�L	�5�#8���R��z�����`K���t��AygP�����A��yB�#'M�S�=q<�5�t�N#=�� ��|t�t����tS��r�w,�h"��J��\��.��mW48,:r����[C�":�ڠw��ˤ����Z?�������DIx�j�s�Fk)ec)��!#�矂f�e����ؐ :�7�&��l3� ����	D՜����~��x��`������BM��	�A��]���&�R��l�Q�ZD��G̅�,V�
�5Ͷ�"�&�����F�-�4���Țm�&����6�\z�Y��8������WF�y�×�����٤3J@��g5��ne��ʧZ@B'=֙��(��QÆ=���u"��ƫe��0����t�pt�����(�wL2Z�B@#��}�ݯ���HЫQ���Y�k�g%��Ǹ_l,�p<~�q���s�U��	�����<��k��9�J�7a��%�ԉo���y,��v�*&�?d���\͗�o�~�b?g�}d�џ�S���X����M��p"���������4�d��<k�z*q�A[���R1]��h��Ē��F.afG�ec/@Q=�mt�|&�caK��q;������_;�?#m�u��I���*_�U�+�ىPo�<�?��9�
�:Z%Y�G���6��^Kt�) +���/Ol��S"N[ɤ�~h�d=�n���;#ЮB��C���I�����	�|�`/Na�z=�w�s}�#q:F�����d-�F�\�b�����r;�kM���d�� b�B�q�
�hd���ȡ��k��5��]�Z|�F(>� x��+獩���"��꽡ͲZ�Y��:�m �w���-��|J���:xH����rC�p�b�@#���+�2sy����Ȧ2�וAu�"[�y�Hm'��};���� 7����z6-�L�ג�E�V�5Z��,S�-���9���JEF/,�hx�4��6�T�cޜ���z~��j���I�oGNoS���{h�͛q�v�~BW�O���	N5��≡p���Qdw@�?��	��¡�9Ц�PL�u���9{�F�v��k�z����iw8��_�P���5�@Pkհ�����_���(j�����Ԙ��5e�5�np�`�':2{���`�/���fج�NwbĂ�Ưz�����drQzDʆ�����u�B�N�z�d�{�T��9݄jy/��v��F�	��G	`cS�����-Czk�<38jOM!n����RKg8�wZH�J8{>�a�r=��^���ί�i��g�}���k1��Ff(�D�=�kQ����>�;�m�x��k����|\q_���
�*fy��ZDK����R���*i睬��I-n{+�y*� �X5�Z�Ū�����|��Q��34ఠ��0���T��[��P���Y(��Rr&�6�!��m�J��kV�])�f��t���?��n?/���`��I �f�����X.U��_�蹤�O/���ʻ�����X��¢ʚ܊��E���*�ApZ���<&�
��9����ƻ_:��6��P=�"���OD|�}�8&3���VT�x}�>a�}�ԑW_�7� }��]�kP��T�,�_�$��J��)���>��Ĕ�����f �r�:N�������gf�m,�&�h$�y���AM�% [!t��b�hz���$�9U\S�Hַ��7�©�����!���m��fs�%���}�n��:�ǖ𲃃߾���Yd�X��݃�A����I5�c��Қ� ���`�y-�vG_�F�^m����q`���U#&#�>0�λkK�����tGP��_�@�'"`�w�	2�d`�NBv���e�����,%�q��+A]��X8��tҗ�a0�r�	FU'����� ���K��%N�A���B;��w8Y\��u���ZB	CBl�Bi�T}��4����!n��!GF> $J�v9�v
����?Ɨ��qF��j���_��CwW�zl6���ԛr�@ 'L'gY���?3��O ��`��*��r�� ��W6%;�VzO��~�+/oP���1z$�}B��'ȵ��%Xc���@τZ��;Y�Di���ݮ[^�cQ�SYv�/ݰu��.�V"P�V�!�Vˆ��h����]�MM?�%uN(e�.�,��l���[�4q�+�oON/�] 0�޹�f�
�x�V������i�ow�Tp�Y�#@N��Ax)���.6�!Њ�;X󶁷�}i6��XeH��#�D)�}��V��k�Sⅅ�D���v�U)��$�����P�c��_A��d�,FQ��E�5����&�K:��s�g�&Q�}�da�aay& a/� YO���F@�$�I�&�#c�Cy��&�Z�u�x�Ƹh��~����/�1+2���%�Gx�%_z
ՉJ���`*
}���G��n3�,��$}�~�n�n�Y��ӵƷ�G<&M[XU�S`�:)c��H��#�_����fd��|ڝڷ�'2�;�\,�jP��� ����0����:�
/�dGGZ�!�q!׋�&)G[q�9)R;<��SNb�ኇ�1����o��>E�&!�֡��ޱTc��F�I������s6�s��R�<9Ҽ�Gc���	����bU4�/F���1��V�.��~m]p?��������� ��"�,sٗ��F;�QBF�=a^Z ����P!S�T-'�f�8����A1݇�$*�Vf06C��M�ƒ�do�A��R��W���fc�3�> �m�wq&�\��e�N<p |n Ӏ ��3�:�f����r�"ڽH�0n�;�$
@�
v;�Ku�H���j=���-��_�ç���F%˞�7\�PQ5-���!�n�"��?�?*�ҷ�-������P����_����Tu�,��?E*}�5��V�.�p�#v9"���3�%��	�R
���'@�Dޙ�����M7�T�o�X)�Z`�����ܞ) ��HX���)�/� ���i��jʨTt����f��e�?@���~�هIo'�)l�(��..y�1�yǔb���_�]w��{{�[]�t��4����N���K&bȓ���� ��]_!n�u@7��s��eW
 �V�E�ǆ��_�;�ӏ�����HR�H�c��/u%���!�b�)����=������:�F���YO��9~:��� !{L�$��O����Wڨ�F��v5��'p�a��;�m�!�
z^�"PH�G}������k5�U�FU��[�%�8�H����o�2��8�uиa-��f�.*	u����X��j�]q��7С�!�,���η�!�=}�����2����qK5���6���;�;���d�: ǝ����:��/s�en��u]���S1�F�Ě�b0p�Y�R�e
�/H)! 6�L�%L#�ч[d81p�[��~i��@��h��)�x�M�~��}t��V/J��eS���lޔ�p�����DT��"�Y��$��2dٗ�l��׎��LT�e�g�H�_�����a큏��I��$�?Y�� �Q"����HȍJ�F���QɅ������,$��򇕑��Ɇ�Z��kl�>��HUyW�Ң/�:4��&L<�������6&:���<&�<B�;����P���Ϩ�B_li��E�K:*t6��e��n����8�f8�b��Í=��j���4�^$]�����	;�=oL� rp?��L]q��L�<
��;k�j�=�p6dk��{�2�gS1�����>Nr��7�#��ןBR&��Rm��tc`<���Ȕ/4C�U��"���X&J�O������o�U��;���]��%�;�r�!�YC�/�U�H#n�'�+W�k�j	�'lO���1)(㽸���<cFZ#�!���lϔ:�F���cJ�PqE�:✯@B�man��R�+�"�E���9�/�0؆��� [��l��w��R×����:������ ف�s���m� ؑ�����0�H Y�h�!k	���*w|Qу���K҉��f�t�﮿�@)8��q��+�r��j	���Ie��)�ۡ�LX>up�ك�xC���q����k:��bZ'��p�Ƌ�A �D_������y��k;�|�f�h.�9��6.�s���zl�p{�1�GR-���v��h�H4����ґ&��o� �����2��0u��6�rHI�Q[og�*6,N�Q 4�$K�x�&���;(_@-T��ӎ�Oy�{9��h
� �)s'�NR}M�jiCxC���G�R$�pe7�G�e`ŉ��B	{z:�q@T?,�58�;�U K�R�$fd��Ԯ&4�ǉ����p��#�f���(ӷthA���[���-W��p����j�� ���0b���+��B<9�D e�;MMdL|Z�໽(��-h�x�H��^�j��2���>#4/��u>�����R�/����=N''%D<A��pM^���z �`n����o���ete��4����DRX_�v6�é�IJ�����ƳnC�_�#Ƞ��M�7
Oړ�Z�f%�3����5��nӰ��rk����,Ɩ<+4�? s_�C����%����+�y��P� �޿~�V��S�N}�̩
Y��S�RQBNÅQ�>�����h���g�d���D�Z�� ��X��U�D9 E�j���r���	��!fA	)�������Zqwh�n3�ސe�jû����G�ztp�CLA���r;�ѳ���6��<P$�9h�L��[��/��o���fj�� ��ɻ��#q$j���2Dv�Ԕ�
�O��<]��}�s����օ��T�����mD+�lha
���n�S-iUuzOjK:$��B�B����>��8��%���PZUI��绛i7����i��\+|����1���^����q�<����������x�͛J��
�������+u���p�� �V�T�SBCu�x4U�/U���|��5aF�xw_��;��=Q���f!T<����%o@fU�+��~ ,�2������w�L|����{��0����/Y͚pjܫ6�+��c�&���=2<&Z� ��� >8Х�sa��3~��7}�pV��&��m�g�^�-KG鐱������,(W�d�f����n�������$!�SF!��hNڽb��t�72М��p<��[L�����ca;O'�S]�Z��$Zi���:ӇϽmv�M�}�,/`�|̠.�@�n�U~�����h���[.�}���>��M;!��ܪ�sQ�i�����P�?u���Ӿ�̴��������:vE���z���͌UU5���GN���l���;`"���Hٟ6���űY8:�wA���]'�Z�����o*S�i@�vv�ȎԬ�_��G����D-��)���R.�3���e�����X���l�Ӗ4�\QWʁKK�Gv��)sR����Г�)�{Y�K�~ӊaշ��=�n�σajJ]���k-��&Q��H6ĩ�ݴ���5<N�lA��OH�6��kJ�]c�W�@��x����H�f�'R�ǖ�9�!:�0�o�MN���$���``�@�D�ξ
���T�y�ogϝ,x�q�d�$Md��w[M� cL�NO�g�(:�唛���L��13��,_	���Z�-l�����@2\��p�&�+�&�2u�J_��u6��9\۽�u�|]Ľ'6�H-�E��&�mf��y�:� ���z�,g�se� {��
�.f\؎MD&{��߇٬	�M�X�Q=U�Ho���.Ąͻ�
	���s;�nB�?a�L��5�����4����/>�K�7��}�������a]T�_�+���5�)qB#�w=��?�-~3�k������5iz�*Бj��fVc~�bI�X\����2��&a_�Eq�er�d�Gͮ����=j��r{+�'��<��{�n�з:��7�6T��i�9��L��Y(GTw��8���E�i�q��i�'2kKLV����������+sP=5�M����.�M�Oږ�yKQxJ�P*b��(��qR�׈�2�Oe��pe�CM�r��fx�֨��N���@������2�7u�%o������=`���$6���"��}� JHFҲ0}j��6L��(�n��S�`u���8���
�M���@�(�4.G u�
��)�+b���b��j^���I��)�X���.��i�FD7]Fڝ�X'n�2�!�d��/���	�N��d��XD�3��l!׾�ۻ�m��Ś � "^�9�5N«���C�xVט�y� ��o¤##�b��Ò��8|�À�!��m��rq�vW��g�{�
j��=Ӱ��uk�@o����[k v�r����5���9h��>�4�����z�#>�S�8�3|��G2Q���A)y
&�!Α���T~���o�aC�\MH,�]��Oߡ88y�������`uL��bAw���sY�����9���ԝ�2���od��^~�"j˖��9`m�(7c���t�/��:��tbl�/eU\,��N��Z}��y�R$z���ג��Pi^��U�禤I)w#�˽�!�[�Vh	�Z%=^i;�D6�d����e�Wr��VQ�R=?���]�M^kr�='�	�<븡�Jcm�r;P?ry@�	/bB�vo)����"!�0�t8�=l��gaS���Y`���NLT6�n9�j��Cb5��@VU���zA�� �){�J��u� �Մ�'�
�%��p��@I���1{�*x�J��6�Jɟ��>�c�o*w���S 	Ӥ���B�K�Y<�|�fN�D�����0��Ǉ����۫w`sXFy�tӈ��)��5ښ�
XJ��*zۖ�%}%���{��UB#��m�[�s�O����)��keDڴ���B����ה{E%g`h�oڀ?x� Q�^C��ȿ4&���0�k3�ةxB��&+mN���DCs�+!��G�մT|X����.�ڞL>8*F��|�?#���q��G!2m�����,_T���b��SjtaP`������^�ʛ��R
7����h�
�%~��0:�g�Z���ӷ�l� �/�W���&�i�d�;��Z�֣��V'�G�7��_Ϟy	�L����\��w�ӱK}#�)��5@C�#�3;ycT�o�����_�:ё71��#F���+
���B>�tON�������M-m8�Jk�=7f�g�`?���TX�Og�d:O�ߥ
\3��\�6V�+�z��{irn��"��ʞc��R��v�y����`r����K�4p��yQ��Z���Qȳ�C����HXL���t­�~��T��J�~�i�l�t�h�N�r�jo�����`z���
�k�Ȧ�B�QN���-5��*N���7��Ve���*&k�	iᰲ�2�Rg�`�M�U5yr&�����j��a<\վ��o���p��z_�������s䶻�@Q�]��x��c2r�~+Z*��k�Hl�2�]0ji�4S���{v4+b��Ն�W_QF*v�Eބ�� �����Ya�O�%���w�7���u�cW����:�������j��]J>�,?�D�j�2]�5��l�J��qx�qz�@���C��=���H�>��x�~��Po �:��Vf�4Y���gz�ܦ^�kK�Jy�!l�d:� ���A �x`gUMRYPhp������t���A�nTN�~1�lb���n����I��� ���h"�â1�n-� ƽ��d�-ݡg{�N/+�JV��)���U�kgz��a	k=ˣ���gV��!�M��	G��݃�D���� '�/��$Jx�b�T!�gL��mz�qÑ;�u{���h�����  ��	CgH��_�5V�O��-H�U���0ғ��TDU��8� m;�L�U)#�|��rimRî�S��)gn~��81�t
'm�XV(6VV�OF9H�n��=�M���v�����;'�i�oV�Y{�2�rx������`c�pG�����^��K��+�e:[;n�T@����n�T��	���I�&3��9�QeGQ�j+7�Y��<�u�fR�Ǧ����d�	�J+�W��j��S��	���z4T:�3����ۇ3 19t=�쫩X��Q�@�f,���2�f�7�KB�"|7
�H0���@��w%z�w+ZԷ'��]=Aw��Y�0+�m}n������JK&Hi3(hEd�Hp�>��#���Ѧ��"-�F��5��!��
g�y&��A�:;���|��������UE��g~�g^l{����9�����Y�b6��f-��c-K��=?:��Z(ͦ`�kLs��/���1�q�/p�6�;��8��=��ڃ�!4����Y�_,2ȵ�a��`��]�A��>e���lj{S��a��CG�����@uv�������@ɷ�D�e".�Hp!���K����NI�;~�pg�A�jA8�a�28Y@�ޅ[�"����rF/C�:��nPg�)*'���ΛVY�+ʄ2L9M�����<�9a�3���Ϊ�uʧ�
Jѧ>}�g)�:i���v9j�F�'�w�^��;��q�(N3��Uk���
����-Җv^�f�0`Mw�
W�#�jBY8}U0.�΅�p�9�#�xJG2R{gx�i^o�Mp�s�Ag�Уw�cq0h�{�f��5Nn��A�,�:2�C�&v��n*H�I�o�����qU�,O Sc�d��6��&O�#@�.��䨝�~�������Jܛ
��k31f�!��%B�y�����TVQ�8Dǝ����y'3ݪ�OP���1��ĬQ�ݼ8&��Ғo�蠂����}-.�_}����yk�؍b�bI5l�bG�̙p����t��?��%,a��6Jo���yN�8��t����� E��1:�Y1�'��������L*�J����δ͝��>&y�.��mF��o%�����O��)�]�I��G��?�3��iuI�Rk�(���+ez�W�AN��\U9e���0]V��e�ɚhS��W ��̊�S�|����3�{�\�����L�r�Ɍ��i��>l�qwY��Z��u��S�A�%i� 4r�9h��|Qnn�I!��v4�2��q�����Jp}-�0��K����%�}�y�Y6�+�p�6��@�3�3�K�n([V�`��)�
�t$L�U�+��#��sܧ\���fm���7�e+?{O��&~�Rö?�E��?��8��3�?���5���|4Um���/�6��o����fR}e�[_lc+��f�C|�����Q�>���]��+�'��Χ��DH��� i�h�@�����#$�I��o �j�����Fm�4�)��x��f$���h��=�;e��z��Y�U������ �v�B�-Y"/���b�a`�{=��8���"���_K�=�,W�`�AKq�Zez���\�t��r�>2w&����XT�S�~��^%\��CWC:�u�Pj��3؎*�O�c҉Li�"����PY�h�hق��zF)x?s덷,qʳc���A^p���2P/e��{�C{���"!{@�a��H	���6�-8b�Hx���u�#��yՍ>K��՚%�?�_y�;Ej���W��7�������e�]�8S�0���
&{�Q���[�4͚��L�*N鎘��]?/�\�)��|(�%��$H[�U�ꀷ��~�u�NE����X7 �h�w�+>1*����DE�	�#*��p�WU��U�*i�#g}�"Ȃ��ދ&+���l��\چ�g�~��'Xg���7�{��j��K<;I >|�KR�n��K�6�M���t;㙘������>�1�@{�-a��r����Zc3����!�+lT{�N�$RǤmѢ�ddD��y�'�'������Dl?2�e�H�s��'0{< W���8��d���[��.˪���;t�zˤ8�s����t*K��]v�d���&dbd*��4��坠?^%�U��Ԉ��M�'j�Aoܫ���
R�Do�sA�!�&*�?Q�ؙ	ތb���b�t!c.��jx{:w�<)�k�uj�k�&�����R2S���7�i*�N6K�ٙ�Mn�����X��s� $��%z��}�D�S�Y0j3�%.��8o������Y�
��R�zn�@��:�J�"��'˴�!����"���D��
��ӽјyv�G�z���i7J��	�A��)(|���X�Avw������b� ��n������+h�P����J�L�J�N:Y�c$*�)W����0Y��I.;]�&��k_��p��5:=�>��1�tv!�:���T���C�s�����=��@��"y�����x}�
r�� 0@�[�_�1����$x���b
��SKF��*!-�G'�: B ���9|m�L�f��'��6���S@e��Хjƾv��|��A�/�L�n@�M������
�#IYC����11Xs�ob�=#�}̫��PJb#|��m0�g8�m�����&�¥�:�T��`���T����̀AiGB�?φ�O��D� ���۸�7cS���F�\J�}��*�"`ę�;��K����������x��������� ?5��-��$�;�O�Ƴ9y`��'��cv�17�)�Z�ջ��8'���F��2Ż\�\�q����:"�z_�������&��/������J�M�'�o�ċ �ԡi������(��������L<NFa���{M�j��X1��<�1;�Y%.9���=U���j��`ڮ���} !�j��v$��p���:h�%l�nY�]@���C������cx^ӏ܂��W%U��)�6��䭦���e��2�$[�K�s�Q�����c����A3�{��l�C��%=9ЬV�@�>YW���a<�-!��� 
�He1��犹��&j=M�:�=�P����Yo^� #{"��q����~�o���Ō�~V_����X�j���tl�/�&)Î��&{q��Ϋ�fo�E�a���t�t,tJ�ae���v`��\"�X4�N�w1��C���cR1-�.24�^��ȕ�kr�������˂փ�Z���?�d����
�����-��}����L��.�i��5n�X����`�{��CU\vW0f%)E͛�e �z�=�̙���=M�[;OF*>q�<���a�2��3
�g{^8Ѱ�v�6�� �d+�~��a�	�����8�!J�����W ���v�Z����NJ��-�h���o��z0[�n�A����Y�hYYh�. ϵ�>����2N�̯�1���zoj!B��3�2^\?2�%��ש����.�r���6f]>�~[�+�XBh`��t*��X�W���O�J�A��-���\!1Y�!aM/�'��ύ���V6�����H��`CO�v�)N��]�9úڙF������<�� pz��p�&����Ƃ����%�/Z�:B�5�W�Ғ,Y2�cg&1��9f���=�O�`��5�I��W˒Wy�_`���s��w�(�F[�~)��8(��;:a��������G�Q*R�t@IlY�8�n(���Ơ����6E����ʑ��]����n�����W0�
h�H�P던ٮ/�+t����]D��;%�.�Z��D�������jt�6^��;T�[���2�׶[����5k�kUŨ>*�b'�)t���چ����ai��n��(�k	��q 	�X��!����W7_�ܜa��<6"3"���3��F7��T�Tn�Ak��;�	�'Vv��/pXs�w�ȫr��p�:m��k�A	+��9���.,L�ݲ������\�[��v2Lq�ם2�>cG[z��)�mo�p�2�Oz�������k��exr�aW���)�*`�/�<�{��HLL��i�V� x75���3u������0P�4+U�L�-��<��o�?3�L`��������S����%`��	����.����	�ap���r:�u��8n22��LĢ����� �3���
6�"z����7������:'=ԟ,�ήDȽ=�N�@5=��s�>�Y��'�I{�,�f6+t�+[o�<�)��Ѣ��ݥj��@v��d��W�~O!�ݧʖvb��V_�Zo�<D��� ��V	��z�\���
J�lS
=�?Q3��Ь!�B&G���)oGv#M��ahhz�]5b��l�֋Y�2W\r���|�����"�/c0㣟��I-�����5���O�݆��?#�!�I4Cqdx�}f�j�z�O%L�j]���"	Sǝ���!��'��U�&�J���4���pqU<w��2�{�2
k 6\	��[��̪��BKॹ�;��,�s��r�]n���T�����`{����j����b�*�ʡ=�l��&I��5�%���Á����-i��|��^H�`(�=:v���]�`'Tw�$?�@�oL?[3��49����D�C�dU��yō?�Xn����l�9I�u�6�Җ.O8�$���e)	�\�@�o� \w{���f�I
>�����X��OA��gm�X�͍9Ζ�3��:\f�.fgҿ�����`B=C1\�&��ݏV�$���"E��"�o� 8�"�����tA��#if�>[# ���׆��}_�:��NM��8c�'��L��I���u�:��?�cu��)��T?�� ����Nd{��t��;e�������	1�t�s��+�-��������������78�,⼕�Jzb"���6ۏ�۪�
������k���=-\۴]����B䏷ѭ����l#+��@�P`&�䴇X�z�?x�4�_���V��h�&�s���}�X@ʚ/SKTw�{���Z��D�L�Jh���է-ȃ[&��:L�Nˑ�O|���-���4
4�&#��n��Z\}N�Z@�y�u�3S�����'�;=CQ�(˻��ҥZ�/���m�[�b��k��������8b�G����;r�Wj�x�ᗝ�͡_̢pxR8����̤2j[9�dC1�vۡ�mt��sj�4����O��3��&ӱbko��y<�H0x7x�K6=首B�\{˶��d�q+����V
�`(�o��~�
l�U3���l`[�O�;�������>L�,�7n����{���%�{6�C���VJHD��?��W�v��R���3�N�:ĭ1W��y脏'\9��t��y]�ZR��h6T���]�z��dqg{`0CX�_��X�eĤ�Fh|yU�T,{+��`��ٿ���F�^��f�����{��A��C�q��;P@{	��SMF6��m�jD.�r,Q��O��}��4S�b	bXHhx�?�aB��9�N�:C�/|��/��4��d0�{_�'��K���fO�r�V����gF�s0{�'��Yl.^��ؚ�,; q�~%74Y��F�*�����:5.-Ѥ�s����s|��?ް��
0�z��\�~��bJ��G��ՠ{���*��v�j�/����o�~'-��]�1�/�����1���N����5�9`ִ�Q���~R�ڃbؖ�%/�o��� ���h�0B#ɇ֞F�ݎe�ޒ˿8�<�*u�8(�/;!li(@�����4�s��w�R�1�*AϰgNE�}��	<��
es�y��=�q�_�8�ݗ901�.$i�7"}V��0��2�x��BKY��g�_������Ƃ�n�{7v<���?!Ď�f��D�B��7ό�S�@2�/�Y=��m�C�G�7_��3f�|�şu|��~�s��<sW\v�&��(�$�����7�ߥm��)���%%F��)�쵌{)�-�~'�{���=��r{�=]��"�G�D�c=������3!�cv���ps�*���93?-�'o��a)��r����{����p�86[˵��[b�6�q����#��t���Ӽ����2�Y��'�i����Ҿ1�t6
HM]����5O��en�Sld��b+k18B5YA7�k!���,:*��W�ĥ��ڽ垈D���!6��>�)�|��}U�B7�k�=v�.A�A��lC��p��� ��&���N͘��%�^������-�A����[�3�_��+�h��D}�ʽ
����w�ఊ��]�F�Q��"��Ho�j�8M���wv9۰�ٝ" �ꂢq�aҡ�~�RN�ߥ��*F���O��P���`|�y4
�����E9)��[i��A2$���ۗ[�Uyp���Qb�̬[`c�/�d��YOƑts{�l�7��y���nH4>�Ҽs��%�+.F�R��x���nJ!���܆���&XSB����Z���vO�M5@�rkȦc�f)��ft+D���������aŮ��x��C�Ql��ˬ���l��M���,��"z�~*r�@
S-�(�Xt$.O�������_T
v�
�E]0ʪ��b�sN��ދ�p��`4)�r������Rv�y'N������HVzV�؆�C�o�C���9�{��=?$����` �����ۅiξ���F��l��J�jn3@��o��4���G]Ɨ��D�:J���J��9�Wߒ�?�p�&Ӭ���w��HT�Qi%W]��8���$ߦxY��S`��$��k@�8:����ހZm�i�t�+F0�eD�!���+�ަbBXj?n��.vrՎtF/��u<t�6��0�Ap�%����sզ�����]G�oU[���������%h]F�]1���~��I7鲺eOR1d�ψqP*�٥�4���w"����aV�Y���n6�~�{ĥ��_$oQ$�o��,f
g�jX��3#+м���p���>P��#Dv�[ᕈ�7/�$dً�OR(�/T�	���=�:h��Y�\�d�\�1"G����G�������.�#$5G���e��ܕ��A38�䵙����Z�5��xQ�k��1S�
�I��xf{0m��M�bW���
�����5�̽�w�����BUn��%��ԭ�����uߠ�;��	���U�o1�^��+O,"���QW���6���~5��}Y�������2������D�{L㾃IS�����?O?�9>.����_}������OJ�=��u?^��i�3��Hl�q���ɻ�L�
��qו�O��FR_q���Xt{�Z�\�?���<DL5�u�3�YP���s�x�o��L}���ʽ�<D@���S�r����ؿ�f`�;J�e�i�
�?e/n�.$t�Vbq5Y^�g�C�շ��O:X&���з��}����"6I�=��T6�w�C�KD@�ҷ�RYN�(%&[.�>L�����uB4KD#1H��?�*x2h�5��7�5KH"�g�ʅ���*l�|�\�
��)L}�"����%[Z��I��`���ց�����o�;Ța�_d��h�x�6��N�o��1g��:;���of��'�`! l/R�ĒA���9y�ĒK������Bĉ�s���hd��Ա��B@(R�s���T�N	�
.t �c@'2���;�fd�oE ��Dc���'L�D)p�X��]�����O�N��Ab Ckyo<h�,C�ݦ#�
ñ$���
'�T��X�&}aCOQQ�I����6��~~{8�T�[i��D>'9Y�J��[���wgμ�j�����v�,V�t�f��5O��]�L�hA�������tZ��j%�����-�U�Ċ�O?�X���q�/�����{�]j9X�p!+zg�Ej&��2���d���u����-[��m��z<%,�6݋[ԬY�W�*F��I�z������Csu,J�ɑ��yW���^�gBz�n�� �D���{��!������ATT	�R:��Hw7H7C�
R�Jw]J���!9t�{����>�~Թ��}�^{�}�=7~�	�j�oC3f�i81 �H���W�#��cV���7��?�!v�ŧ�=J4N�VOh{���	��DjT�N���Rd���b$���J�J=�XC��I��=�G�X�d�r�:EL�& ��$)����,�*A�k��6�����/M��]4� �yuǀ��#�5Rt�CiE�Ѓ�U�6��i>-?o�m:�!tU_���A�=N�5��(�ME��!Uh�A6�]�[���J���ƹC�X����^5��Ĳ��-� z�3�z?��T��8�c-w��E�����ط*�&S��R�������S:��_ ���ƴ��+���؂'pU�`D��p@��hקּ[!{�p��"tu��f�MT�-��D�9������t顸�o�����Nge�飯�e���zrݡq��A4/�1ʣ0���p5��t���G�8��Dȶ���L��u���X�8�ẽ���%j{q� :���l&�.l,�<5ta{���$˟�{����5@l�ʪ����{��hX���Jo#"XA}kh6l�L��q5�tn���s����*%���{0�u �����k^+2����M�R"w�*/M�$��:����ޓ������[���*���=��!��� �"�Nʴ;AJ�2cǋ�LG���웗�xth�AOmΙ�o�K@�e�k��IZ9�-	��|�)t���H�I���.�����θ�\�{I�8�J_��5J�����ا�g��G�w���I|�5:M���)��Aj�ġX�z�3�c�[��+nƲ�ܩ�k��R�N��a�r�HrS ś-%t����.c�
w]�`�G���Ӡ�b�i����&��0��a��\�U��� �V��K5�3 Oj<���=���Ņ��tm�g�܀�ȣz�����s�_�,����*"����d�/X3!#�<-׼&���m��� 88����VMJ5,վ�`�����em�����;���z�~;�z�$k݉��;/!�����]T��TI��%����&�\�ڢ�����SCbp�(v@�l����:o�͟�V�I�u����]л�����!����?�a�<�'��p����ޱv{g�⵵2dM!f��� ks��6�t^��^U�)�����4bg���>���&���w�ݣ-(�q�m�:`C'�<�t1t�9�-O���M�I�AX!VS-,��r^q��RzwO��x����1
Թ
�ߕ��%�T���/�<R�?|�H����o�q!2������9P��T:YQ^;s���/�Ї^���Hrx�ݿ��.� 9$P�
gp���T�]�P��H
�,6f�����i�UH��he:͂tBhe�3NCZ�I3(-�:24���!:�QD��M"�xԥ�^/.�6�LT�&8)Q�+6y����J��o/ �'��>g�jd*d;���y��*[�h�(�z`n6�{[�P�J�'�ښ�V�|��!��������(e��eҶ(���r����o�Az��q�+�]w�Gu/��x@���T��B��5(�g4����ᦦt�׼������s�4( ��U�W�P���(���F��f(���?Z����b�"y�\ƨ��E���Q���Jd�V����k��]��� �?��>bX����le;fM���̥�G:�O��.��rH`b�s���%t����5W���r#�_N6?2U�`G=*�8���,����B�H}�Lb�.�Π��~i�O,7h�`)��o�o���^��8$H{�q��a�4.���;,QҾY�vl��ŻJj��J>M���^��2+R��c�>�B�E�0SA�2V�~�΄q[�@�l�TJ�k�����*o΂w��4i��
w��9�.�!Ζ���ܵ�	?Giv��o�&��F��Z@7�	��&8�l�c\T�+�?��������L�"�X������23:����m3J^���6��\�s�%X�Q��޸/v����ib�;n� RHu'uµ�r~�r���Ͼ�-�}�L⌲K�{Wm��0�/�ڃ�V�j�(�o��w�=}��=�o���e�Vn){�Jx� H�=�8"J]��՚'�v-�����l��r7%ݎ��5���P���W�����6�����2Z<��	��w���L�?�+�	��_=r��L=���@[-m�Ŗ���Mo���_�S��Oᕭ�A�Qu�t����K���z�>�ѵ��y_o�bR62�������%�xj.��Q���a���eB�민�]�����^�kMoן�/���-�9��:�侮=7<�J&��OY�0��-���/���-�@(��m�B�ᣝj1�fk�=������s^LT�o�`�H�A!���)��	����Wo�+����)����jI_���tR�7�Y:=h �`���U�=���'�6/]�-�Sd_���r�#���H��<5b��W��R����C�^&�~-�p1f�o��������?�`0g��?�<�����$�Q���6��؞X9I�������2_��	��0�dD֘�]���7�D�%X�/5�5ܧ
��ރ�;��D,�K�w]d��c�-0��9Gm��H���݋�ͭ3D�-z��f�����xy���_�*��E��80Z�V�e�ܑ��1�-�6C��'�����J��?��\3�f/:���%D�^\>ޏ��#���)�����?��`�e�Ѹge~�ypt�3�6G�1k��

ñ}9�o��4ǰ�hP����`��p�$	K�S���*���ڛ����b�~>��(\u�!²�QMB%��<L���:H�>��h�~�(:��N��-���M�x� I��|�g����.�j�,,�w��;��ɾ@��]�=�#ԥ\�y�v4+�b7ER�˲jaڲ�Z>�y[�Y�n������]Mu�U;H��$��P�#T+�O�˱Y��}ek�(��%R�O~��k6vڛ\�z���Q� ��>�f0�Mݟֿ��ٔ���M+��d��W�~>�����~s��'q�'��V� ]��;�9y6��7Θ��6�9�.	~Lr���Atu�_����P_����� v�.<�E�Ǵ��������ƕ5��4�]4�y�����+�ɖv�QUɣb�g����H�qh�!mãp�;8�|捔W�RK�#�^����; ,��<����n1���-�����6&�z���۬X!�Ş6�>��A�r,���x��7h߾�{��{;QKA~��}R�Ӣ�}}�7d�~B��� }���ϣg��:A7�{p�������������w�y����M��
�ʎG�꺣��!�Ş6$��6�5:�DV�	���5����^��O��R4�_r���m �x���]� �����y�������:n��	U��j͒ʖn�'�͖�)0}Fq�U�I��\jBf���#]B�G?�t�63���{ϼMg$Ĳ?"�ر�&V�# S">-`GX9�\���f+M��9�+�_� ��4p�PňPw�@�K��b�|�Z)�ƅ����a:��	rbӯY��ո����4(K��:�z&��u���ݟ�Y�J�iy�ۯ�Qc��;��#�XaH3��ł%��zu�(�{f�l���ˑ`�׍֚�`tٍ2 ��>Xߵ�_��@��׺�j����肥�<@� �t�&ߙ֒I���Uͤ@�]�μ�p����L�yy�D��f���I�e���c��R:e���4j�Wia��S��ԵV^o:�۳u5H�|�[�,��,���-s���Ȭ~���~�E	���
Td�MLcj����S�|���i�o�C��7����V���}���}��p�X����E"f��O��~��������e6xA(}�¶@Y������XI�/-?Շ�.?�f"~)(׿�V���8}\��PU�(E��eǠ5>�38<��I����
���[�5m�Oט�g]n�<6o8�oq����]t����%y��D�(J8�%�{],�X�u-%s�I��A�����2Y'�/74���C���(?��t��I&>���2-�ĩj��{E�{L���<o��菙WMx��{��e��S������=9ՂX̏X!K���Z�1��Fqa��ه%}�h�� )�=�7��d疏�*)�T�]\�GQ+j��cQ2l�>x9d��T/%܁��lձ�����o䷘�E������s���Y�(�ò��l��X|ak/^�)��B͍����an����!�Z�>h@��dw��F^#�+�~�����\�n����o��g�Gٺ�$'9��K0A��t�� ��ujVhPns��py[ӌv�9�p�<�W�:�3~�����C=^�ogk�"�� ��I�C�H��U�n�QA��j!t�H�Ǣ0=G��x�O��'<`����d��'"5(T�6���Kn�5�J4��t��^�7[������.���
P0�E�ﯤY�?.^����7O1��t�*���a/�1@�j�f�hԚx'�Fg����a �A�&�,�7�r��"9����?����I�tH���H�TX��d�w�M���G+���҇^n�ALbȶl�V=m!�;�AƢ������>{k�H��<(�e�߳��G���f�j���k�\�aU�xaؑ�j�$!��n�a�oĩ�|ޙ��7(/1P`�#�	^p䏄<��'�͉���ﴔ:�Y�>(Λ}�VXUc�JȎ���g5��m���>	u�;3�/������I�jf�xؐ�l�L�)��F+��O�x���y�|J+��%)�(���G��7��)�K4G�*��lͳ�p��g߆�ɛ	��w�x-76轷BTr4n[#��M����PF=�b�������@_����@}������iH�M6�d��U�P5cɓ1+# �J�:T��o����v�k�����oWwj��!TǊ%R�1K�m�{�񝻒~3e�]���Gc�~�k^)]70�~�d�Ԝ"\Q��u�3 P�+��k�o�/|p}�:ݝ�l8����ک7��a4�Ԑ#��_����`rOfN�;p;�A�R�觔	w�qt��ʽw���� ���ͣ�/M����	K�����V?{D���&	Pa�����W�஀l��`^��E��G՛]�Mp�!_v_E�Z�����_$Y�e�L,X���D�RT������Ь���2���O?��Q���^�:hɣ�RAGq�gq���[ET��Z*�a���O�g���� ��Ǫe�~��Meu#8�~�����f+Y\iH��m�,��d8H��:�D>b���X���UHQ���޻vX��QV� C���w}�xD�b�%�n<��DJ�PYd��0<�g�J��K�C�oA�����D�3n�C8�����x �|f�qE��SUr�% �N�{�1`V�W�]~�%@^�F7l8�IR;bV���l�v��~����wv�����6'�Jߎ��>�{��^܅�$E�7H��ͣ4L�C����1�&&/Z�������/�`^֭mC��;�t<~kH=B�۝���;�{k{ё��@{��*L0��'�uw�k��{����º}*<���4���p@ZhR[M�U	���L��	
e��j�����$����4ɜ���;��������*5f�煫b��ªx�G/MƊ?ho���0� w�;�_�&��Y��7�jP��Zm��e�D��,��G�Ga]���в��b,��y	�U���ü����%}l�I}MA���~0�=�	S[)L(�z9�wjc�6 ��}��'�*f��P5�.Rظ�dvM<~V�PiP~%!M_m�w�X1���|���W_��	��D�<{~hG\�#��m%�Pnm�!rl6���dƊ�ؓ�֞ow�zVYa�A���ث���D�V"���d�H�OGq�G�a-����F�Lڠǫ����r���]�����7H�*��f�w�F���+���"������n�W)Qm?�a�{Ǽ�B�֜�[w���),\��+��"vO��c#�Q�{�b��"����jl����;����������iI�9_G�X��K�Bgtt�ݡ�yYUGe,��|.,n��֢��
g����r�ܜr��r�^+eԓ���;�c��T=�.�dR.����zK箕���v���竄U	S�N��4������2m��S��N��׃��-x�=X���_ ��h��s��� Ds=�7E\k�d�9߭\���# u�le>�͕�ſv�*w̋Ö"V2�$l5��^�^�Sgl�[�s��N�h�R��tn3��h&?�����>��o=a�.�^��\�f��ż��ݨ���q����D�9��;c�F'�t��Fv�qa?.�+����j�D=���is�����UZw��n~�i�PxE��gz`��;nU3|y��$�����E����=����jʄ��t�k�|$X�e8�c%#�X�����Ht�G�ol�@դL�Q�
%*)C������Q����+�`�pKT/r�b�������bP����3�-���/ZO	�@-P�->i�Ns�Z(}
�?���zb��Ј����0rP�.V�ro���*��z(������+I�xJ^������>���0�[Y�^��=�����_3x�Di����������T��q!�|�J;�]dY~eg����)�i��QO������r%��?�N}��5�GJ!k�FƂ?�Mf8n�`H�j.>XB�����f;Q�� (K}s�YP���]�M�	`/����������w�>��O��'�����mz$�J6�G���k�C�Ϙ��cP����g ���N�^$W��QA�,u�f�����O(}G��&}����v���=?�|��Z�N�W�%�����{��2b O���bc���'Р74DN\4gk0��>����O�Z̭C �� �sd�jP�[�q�CAM�2-�S�9�k��������)�ּ	Z��Y��_�bg؆l������Щ��Ic�%����"�@I,�  ���.m�Ͻ�q�rlAG:M�N`�?#�R4G���CY7�৘���l����:n�0K� BW�^}��'�D���t��spR�0|l=tDXz��Ǳ.��c�>��.�Nl����=f;��v.|0����O��?,�=GM��z�x ����������[^�^f��Bd�)��巉�ER���#�w�.�m_�#sj�a�x����Ve�U��x�x]Ȟ�7�^eװoH��KC{�^�q��v�~��Br���5/���R��%��� �ǹ����W��������cn��}&F�2К�-lʴ�
LN�H,���g>�q��_�
.��oS��
�Ᾱ�ϙ�p��&d��I�^�Soh��Ɵh^LU%��by�:������*��`���j*IS��#-ٴ ��P�h�ʂ7�u�����ok r�i��σG�n?ol��nj���l�γ�/��H;?�U�G���?V.��g��|�j�_:��CҠ aњ#�#��9�
k\�eC_D{��d����,��ok�-��GG�zG^f�����w�1mPe,1L�tK��u��|764�MF���@��OGIe�Wj���3!�0�;�g���}å(m��A�7%���s-*���6~7���%~R�< =T�s�`F�sEgo��_�n����'�ִ�o>%�0�Y��tj,��A�~`зn�TFY\קQW1l�pz�l�4r�"]�/��a�\P�'c�A�fr�OPڂu�'H��.�5{oH�B7���������>���4���C%ƪ�a��@��=�����s�"!J��i*�D����3/�("��)��o`9EF%�m.�m!]`��H��웲[��VO�/P�,���~s��Q[��\��ocߴ������eHO��.|8dA��M���Mu5TG-�]�bmf��>8_Tr�C4c�
Y6.�4yz\�I�Z>~�g&��&�0�k�	�x��M������&'��ٙ(���_���� ;���L�;C�$��������aj荪K�	��m� �N{���O����7�ǣ����/�=���L�FP�J�����.A����R���]�B��j�g�+�#N�����O�fOp���xO�Y������OU�E3Y�!^^���k@���٬�5��}�Rme�\��{z�k�j�$7\��;D���Y~<Ll��{}k�X�p�U�DB�Pwh�ta�u���O�����²�����B3k�$���kȂ[3��`�m�� \`�-Q7HgA�diw{:�GMf`�W��GF�.���
�u%.�R�m	&��T�͠�������� <���[W]l��=8�s	�5<8qt@4U��Y���D���J�����������(��'�&�!BҍM��{��v���f�tb����e
� $}�NL���� �\�����Ypۜ�7�N��r��W@D�+�t$\�OI��;���E���
���	M���lA]�]�\�W����J��}B�p�L�П�>12�c�A���E�8�MT�2$�7(��o
��E��U=���J�$��Z����Q��t��}@���4�ɻ�+�_���6��I�����I��ųDa֒����<q���'�����{c�K��}2���ᡡx�t�M7d?��Y>��%��F�%G	h��kh�(�����T~�4�z��b��)h�_�ߒ�h�Я�q%�=���{���i{�FA�7�"������V�X�s�r/����$;�]��L���}��9�K����Sߋ�qr<�6�mB���ښ,����	��B��NA�������ѣ�|j�s12�]����v��Q�v�{��p�����A��O����������<��,
|720���X*Г�W����ݭ�%�)�����p���f�q/��}��~����9��I�2�е;�)n0)F0U�a�6�)�Ǿ��&�M�.z�lP��Ļ���e�gS O�!`���N\%c�i�+�������;խ_��b;�Z� �L.��\:�����:����ܰx�ӻ�����,#�V�gZ���l���6����c#)��	���`i>;�-\��Y]:%�Z���W9;�ڲAK`��먳Q�#t��9�&<����-�|G8���r��F��o�3bf-��Da�5B�E�K/<>��!���.�������
YG;��F�9Lo���U��X#\n7:"d�����N ���vOs;ȳn�)�w ��]�p��HԢ�p7H.YK���i�83�������H��[��a���5,G [�G�b���y�6[�3y�2�D9��\mU���3i�߮�&����(��w:����,}Vȇ��R��$�O���=̐&��8�NF�����em�-aչ�؅�
�(�*��������P)�+J<�;c#gb��3ЀZ\�G����:�4i���3)�vd��$ �]��'t9pC�X��8{f����~�hR��o~�zǪ'Dѥx��C򌧾�<�I	�0av9eӏ�M)�|ڦ	���޿Ia�����2B�Ρ�C�w�XW�b�����/���=8a�Z�zd�k]�|�_�^��>�|��/
;���F���"c{���^/0@��o����Y�1�1,
M��]�؁Ң�*��+/Ei��8e֬�%�P����ۓ�+���W��GQ���
�{,1���la�k�1K�,LrU�t0�8�����f�~\�Xb9��0���!��$��tM������3�T�Kj���f�o�,&Nm�=�Y;���5I�we~`��1�X�=�ڣ��B�MVK[Y��f�&��U�K��<�<[�ǜ���zK�"1u�s|�͏��,)��o�mt�/����C5��zU6��D]����Ok&��N�_�Ҟ�&�n�i6�71^y�σu{�X�Qh�_�	(6����l����=a�I�Ez=:�����%l�Iͨb)���,v)Ġ?�.ye��,�d�Ɠ��
��-��QoC6cr���(�,)2~t�7s�m�@��0�TڗO��$�z�0�Ӹ=a�˛ȧC0v�^C��	{�2�+.��*?`��+�m��.�E��歚C�����ֲrA\{#��7t�fLct�2�b�җa6d��{_	��ڛT��K3��?S7{�u7o�e�J�~��-��ß����B�\A^��;�E���R����m?�K:�Z�]YT�C�Q�vz��R�x�XjGœM ���n�O�$��u�oW����ĭrl.���/#�����Vo
��x�)�b�V���^���Д5�gN՗�p{pΈ^�F�%����s��Y���|]�建�0�k�+U��eEn�	&��˻.�HjfH]5U��~����^��+���8#�qq`�1v�Ҏ���C[�h�k��q��<q�����Z��,/�K���g~����5ɢ�c���-���bh��3�ԭ��XгK�=�G֞
�1��Z���h��yyy�L��O9����?�פ'$4�5���q|�i<J�亽+pL�9WCm�F)v-^)���`�`��?�^�ag�n���j&E���vvFEQ����M" ���=u,���x�4�ſ:W�ẘV
S�+����U>Z�-���cy<x0λv�y���9�k����xz�V�j'�VV���R�]��}X�à\
��n�a<�=_j��ܞNU��kˣ��Z6�*b����\�{D�p�\'��!��V���*�ESZG1�LP�c�y,��fh�R�AtB�j�t�ʃ.mo�{��Pc.���J��۞>'ӈ(�QV7���;��F�QU��y��-j���m�~PG�|�>n�kn*�e�#fz�4��LE-�(� ���V�/~��?R�(�Ms�K%����e�L��d`w��Z����/���ݗC���G�O�G��d	���j9դ*"�"~S�.���gv�p>��P%��r{Z=��"���l1��e��ֽ�;+�[��}u�ׇ�x̥�*�0lN}<Y�,�t��Lw�[Uəu�K�>�si۷Ծ�^�̻��#�UC
��9y>V�v���)W���B���e
A�q��H�6����?�Lds��"ڐ�v;Y?*��й�=�|y��U��(��Q����o󋨶�a���\6�IP&`R���5/���_�d���oyA�:^ʆn��Y������^�P����|Qji*+�ɟ���L ��L�Hy/K{?@�{��b��s�~E��f��lJ#�7��\��\
�t24�./����qR������m�E�F���-ѫ^��SOMwI�X�-�`щ��<�pW����LA����?��6 05;�1GU��P����
-L�ܾ����14{N��Sk]7,��s�=�;�1S�Of��WW12�˩�P��o���ƆEmJ�G�|�Aڃ�4T�X05���5�C	4k[p����C5�Ч�r��$8J8�~���H�����L����^���j�YܒO���(�]P6�H��=ef~�������"� ���/�^�����pU�'S��|�C��_X��ܷ�_�æά�$9x]�%���vv~.�y;f�f+<�zy�]xP��)�A��l�R�39�%�	:R��<��&-��alGQ���	��ߞ�W">Աh;L��`S�>Ĉ�w$0���j�#�Bѽo 7���Rr�q#�u�V4���ON��[#�PowS��5�������!}c���ӎ�C���iU��Y��HĆ�C}R��P�	7���7�ӕfɈ�l'P�L4��G�l�o���f��J����Q����K�����U��]g~������ψ���y^K���B�w�w)�s��q�k��M�ĩ�L|���{����κ{S?����ԥb�`����|�و	��Z��|t���;0�X󽱝5�?��P��m������4"�^M^�cc`.���=KN��r��W����O��3$e�i���L{��S�}�;����"���ꃮT~m��	uy%@�b�@��KG�'��#���N��m�'�/�b�$���E��5���y��^��i1\�8�)�$y���� ��IZ��/�Co�Y<���`�����6h���������;��q`����'�|����WH���itF�A}�2���F�M�}�Zhz�@H���v�Q#�\��T����ud��\�k&���*V+���.�<�G�n�x�Cb�;��t�6�P�kXW x=�e?V�@ނ�ꍪ���/H>m	���A�#�ݎذ'_����#��~@v�,0r)�}`w�ķ���S���ݼ�P`��f["��d@e>1R�P��h`��emeM�����,�}om�����T��%mE1�Gߔ�9Ʊ�v��ؚܑ�#pߔ '��V��m�l9?�Pk?Z�.D�R�_]���;�$o���h�4��-p��ޒ�V�m��΋�>�۾n�dgU����x��Sh�$�_��șZf3�R�:��C�5�x�	�k:���L1��kv�4���&���ֹ~k��HVz��\S�(���d���idY�e3e�1x�o�iʒ��վ�_H卌�͸�W�1�y�M��9k�$>m����i� �\��5Y��w�]d�e�I6���;0P�?c(�����zR�kӇ����"�r��FҶ��ʿ��a7�9V'�L�;a���?t���(������j����gPVف�W��q�$92�A�	� ��^8]Y=8&E�k�E0��I�p�}��!����RU`����7�����;G�5�L�U�P�k�.g��K�wK�o��8�, ͑�m������ ��Յ��J�#�X:��p� qVS�����s���2����h�H�O�N��ȯ��U�X�*�������>?��D�(҇����ǅ�1��D���pr�>��ŗ��*���mOA2��.Z�К�Cy�ޟEcB49X��(�Z�HZ�fZ�Ju��f���_6�6H�8��dǠ��ɮ�*�x��8�Ã�eo5Y��M�հ T����r,���8��J��AV���ʜ�H�.#m?$�%�~�4��)'�;H]�t'qCMF��a��*�L?�@���o���T�dʅX��a��S�Ĩ�8�}�����!���5��}�!%B��[D1Ι71���N^My�<��U�V����\�qTL�Ov��Z2��7�g��ݍ-��B~���%���R3���+Y�9??��fe<Es3mZ��'
�������6���C��������V�&��gf����Gm�Zd���4!�b�B�]i_�N8���\��$6���� �1�j&���v���Rr+ܠt%�X�W���ͥ�x�zꕱ�,���T[,����d��9�����¸��w���ކ?�y@1N�7��B��J?$L�Nu��F�H*���LA0��a�j(Q+Q��o��� �}���0ƹ�����)���1����Q���k�2l��	KҮ�̄�Ȼ������u�n�����H��z�0�'�f}@�
rA&��"��*�.b=��./�Ŷ*�V��k˵WPa�l�C
�]�KU')U*A��x�+�6�Y�mI���w�]�L�2B�Deި\#�3ɔn��j��~��ӕ����{v~��҆&}`��ּQ)O�������#T1��C
arn���E���}CP�m=�3)>�h��+��{2bZ�R��C����a��Ո:o�m1[�f����M&*%JT�TRn�~t�쾢��be�Wjf�0��.��y;�'n�w��O�E�F|��ld&�Zʘ��m��R6Z	Ǯv0_���Ft׆g	�u�O�%��3*�|�u�B��<P3F/`��;�'��ƾc����e��8e�F�Íd��~e��T���r�Ԙ����{MN%�T��Q�O���F��v��U�D�>��76�8�����$俯Ҁ����Ŀߣu*�I�R���2V�����aa$�l�_W�?Y~�kޤ<�tW�6K&��yHo��;uv�SQ,Ϫ�Ang�X��3�RC��R�G˰�� �ogK,fm���^L��3�J�E�\��0,�w�'
[(�?؛�*3�Zd~ �l\��r�Rvŋ�Rb��×w�w2��P� ,�!�
c�X��/���D�zc��b���ؙ/��YH�47�
Oɘƨt��^�W!\`����hG��x�Y@"w�M6W��k����e_G8��)-��1L/��c���@Pf�<��V�.E���>�p1?��u��gzr�c"HR3ܬ���`\G�IcX`�X�I�Ӱ Tef���<<́%����cc��I���07�p�>�W=d���\����o;
MO��	��^�m+����Ll�������A1 ��B'�9��.K��6����3[�*�%��`��~,L�������K�vVh�IO����hF���W��0BX�f�f��gM�p�R!�e|������`"�n�Fж�wZB5»o}�u{]v��I�Q�7�����2���S���D�s��Gv����ɠB��
��f��H���1Q����WܩN;ʁ�(�\���t]��#�Up0��դ�dp��R��5h_\/S1L#H�{�e�)`�ݣ����#Vu��%R:��F5�>!۾��˩��A]@���Ͱٝ]f��tFｈ�5 �ZI�S�`��>�`�E��U���$�jbK��[����Z;�Dd궷��� 1�P�A��pW6�~o�>�W����XzNd�O���H�r'4���������e��+�FH��@���RDNC����Y�Y�i;���5�*�O�d���9ޕ�g
�Y���e<11&4.��7v�7�j�7��*=�5TAkR�[�8E5���'Lob�����n��v�!��� ��c�lyE�@�l���K	��@���G])7E��>|�e9��4t�n�b�=�=a���U�d=R����Q��qR�U�n'jo�R��C��V��^��*�X3��u�Fu��Ah����#t���T�J>�Q,5{�!�½�*8�%?t��)jlG�J�#K{Gь�]f'�{�����x�I����ޤN.˟��UJ�BĢ��h�~v�Э�a��d3&"
�tP���h�L�u&@xn_tW�>���ȅ�d�;�����K�\�f���Je��ߟ.��)FP�X����'L��4_��Dy@�q�C-��w@]�r�r��2�A��Y" k�;�Xز5���;�⤟�5v�?bQֺN�V���Fz5;/�~���γ0�Y$$����s����׷=����o	$���KZA��5+��p�0MZ��N�;_M�\~w����V㋨K���3��,�vț���9�X �V+yOҬE:�e&?���Σ3ϡ⭹+9U2�U����"| �~t���y(Vl9}��W��b�W�;�\�c�ò��U,�ml�B��"ݺ�AD�j+��1�9������g��+��3�c���l����w�2�/%g��^nG"��!N|{[1om�������A9w+ʒ�T��]���ȯr�9I��~��Xh�{$rtjE5�	�? ��J�H���ņz�$w�g���v�*���L"D�V��;����L��(�M�8�l%�&��W]�A�W�Ki��wK�4e��L�ȿok�V���o�Û�eǙq�q�ȝ�ޕE���N}2�` 5Y�M������}kw��gj�a/��,n"����{����2Kl�͝9��fړ�e�$ᆽ�`;.���iIe)�Y��8��գ ��8X�SK���d�!�@���������~�m�0�@��/���d��y?�8iFF��S\/��}�I��^�ު�"&�OA�&�7�O�*	ZdV��eA��p�6l�^��B��I]��O���O�.}�\O)ܭ�t:��Ô<�-or��K�t�A�Ǌ!��Sj�,�G蔓�����KF=f�顈�oy|?��qx�*[�i&+��(*z�T�u�u�T��O��9hF,�T��g>�۟���]:���V�b�h����_����&��떁3�zPᏍG�	��r�wV�1��Օw�4�:Zs�s�v��H�F�B���?{I�,�����m��]:�O=�����l�����r �񘓧#��'ϝ�cz^��f8�P8^]%*\�~U�Z��]	/���ʯ�cPΆB�U~<���"��\�2���<���+��+�K�bm���=��\x,�3���3-�V�V0��6��A�����n�D����j~;x`%gс�?�HA�d�M�/�o��$��*rEW������c��:C]�5=T����3���3��C�Å#�!��f��]�ۆ��rgu8��}ߌ���~NJp�P�����^��Ma�]�W`M�?���Ҟ~�Rb�^�z��X���/�w����T����l�{X|:�<�����(�Ry�;M����h7�.9+F����>�]�歱|��'*�v��I�����I}����94�3��i�d.v�2
��q���	T4�XUĚ�`�f�����2NL���t>�Qk�t0�B�c[���+-I��W�aP�#K󸕭\_��z�@��-7��D�Ǚ��ȞXv����B���y�[\�eZM՛��H�Y�;㫁k����X��t5�:���i�%�]Tӫ̈́<��rߴ�{�~�
7��Q�7�r�т�w��_�B�JĐ�8w���u��x˩J�s���j�q����+�BM���C�?��*�G����oʛ:"se���\��@��r	�f=���e�ۻ����v�V`DeH�ExK��2@[���K���d���Y.��ڥt��ԲVʝ&�ј���������ڜ�/OƠ c`]nd�x��fޑ�����y�q���]�o���b'"����B��ގ��ld�$�f�$xS��V�zh1W����(aߵ���Rh�F�Z��ZrGWG���)���#�K0��8
�$�6��wEy)��o�k�(y&x�EU����9���uʻv҃�;���տa؇m��n>�T��a D�i�\��(� ��@iW�u����WD�oƼ?;�+6�N��S�F]�nUW����@s�����O]��'� L2ً���ߦ]�g,�8�o5A���$P�T��Ȑ)z9I�8�l����	���|W�Z
쓧=V�1N�bdF�~��	�����79]Y��T���� $6Ɖ>�LE���g�դ/(W���?Vz�,��P~�=�M~�_�;�9*D n��U��#M���PR:u�≥IO]rV���o�<�z[-�\��&Y/45�,��7�/�(�m�k[{y������Y^�SI�׳��	�]"=�C%�M���s�'ٚ�v R�M�Gu�Vrvƃ���2N,h�E��P|F�\A�t�A��E�}���7j_*P�j��z���9lÛ�Q[Y�Q)�މ�����3�Nj�h*_�/�<�K=�l5l�Z$��z��HL����?�ӂ��S���3^
�*w���7Ģ��z���^����.9,�_�j�C����� ��P;�٨�)���Fׄ�r��Lz���O��2�ݗ�I߹3��fU���r�$陫���z�(��{xXVp�`3*QA@W����3��$IR�HN�$I����4��<���a��}���s]��s�=�������nK����f��'a��pF�{ּ�&f���03rx<�u ��`�oԳ�p���O��z�+)*Δ�>x���Ѵ��W�I �X�g1R}=��9zF=Oi��۷|0�f���|@�iD}�u8� g^0�^OS��`8�HJ�	�������pe�?e�P=��ĺ�����o�h%e�2V��7�$�=꬧�ؙ�>�Y�)��y��H|�*ς�Q����#n�s�hjOE�8�s>[���7�8-_VSX�_�u����65U�16��M�6��f�k݋�j�����"Y�ћ2��_r���Z��5��6�h������,��T~���%�n��(a]U�Tja��f�.�η}f�����T?3æ}�'J�t�� �=<ò*O�Ct�u�Ps:���?8Ѿ��^�ޛv��c�c�	���3e/�>�M/̅����ŉ{�rZ�Z=�Q6sm$vc�5�(`m�2P����1�ٱ� �T{+?�rPm�6}i���)�ĥ_�'\�&�rB��#���o�T9����Ci�����ZފcE�dg�W��sU]qL����a�Ms��@�p* ����k�MWUD�$u���<;7;�ժe�;;�g�vДq�)S������1���E�y�|ѥW�,?��x(�Y���[����|�9��d뛞L�u,�4����tʬ[��ð<N�p�(.��
���I��J�Ȩh��_vM{����3=I��sX��T`P	7��Iˎ�͇<�I�E�����}�S�� X�m���ӉN��]ݿ&����_�5ӡ{4:k�����z�x�5�|8M���:�7v�@�d0��V�ڞ6ۭi%b��G$.�-�Y�Э	�v.9����u�vO���*I�\���,mǪ�1�����(��2���&��G���j�~�	�F��|J�M�9�����l��A	��9�'�����w��,RY4��n�{߶-<���G��z���1���nc$r�Tt�	�9��F�V�5㢰5���_����4m���'H�qŠX�^�.�1�z���gK�I�ǡf 8���׮#����<��ư���P���uQ�Ӳ���'sOm�æ��18�e;	����1(����;k쭛1P�m�دmoi�6�E������8�8�(@��6�V*.q��T#�J����Ǹ�6�_����(7�W����))��q/�%��l��B�������|�s�#�ؚj��蟸ab�$�"�)�������t�*�ܣ���6[[^����o*'%o�k/oׯx������#ʞ�$0ks�Ӡ�IB��66�i̥5���?k��T�����sG�vO����N�����(z}A�R��v{C��O�뱾NУ��^V� ����ņ�t�C�(1�(�4WY�<��cW*
�����6�rQ��qZiz��c;�4��
�מ��� ���ԃ�J�ě�K�@�l|��G0
_�,E�������W��0��
���pm�����`܏C�%�u�镠X����Rps�����t��hVn}l�@��Dg��Ci2[�ffP�~���fl�W��ofҴ�]wRP�r=���|��M�b`���2:��X����_�jr5<���閼���;ZcƊN,|�*L��@~�X�0u2>-��$���ϮF%�i�+�T fm��P�Y�=c��]E�ȷuN0��1|I���f��g�����8�"���μ��</)��ួ�>�[�*�A�Ot<����8���MnFj*D���P3�Bo�������s�X��� r�0��}5�ߢ�xՈW�w��#��j����^�(�]a 6��������e�L��]�FB���E�|��oŜ��	����A�Lo���~��o#3|�QN�i���t�)�+�)�3o��xM\�9��[H�ǉ雂h�E�H��+�=��f�8r�N7$�D�E�(�U��S#�Ds��S�Ⱥ�Քva:��d�S^3���we�V��jC�y�T�n�KWPES�H[*Hې�����68Խ*m�un,�\�SZ� �J��}��pIn�P$⪂rN����C�'Q�Ɏj"�s��Ď,���J�<�b�Z?Vn��5qnU�L�Ꮮ}B�l�]Ĵ������q^pĞ�z>Ɂ�3+2N=�D`.\`$���H��Pp6�9�����Rمe�Q�� �v������?L07��J?�o�Z�������:]�-le�~�Ĕ������yw�R��O�X�{V̯��zy�P�!h�Ʌ�K�� o 7�eڳ�Q��Ƭ��>J�O�4�A�����)��S��9X�f�/ F�H�m�
B��c�l�k�[j�j,�?����oZ�}`����,�H�H�T�u�.J=�J����z���8ORc/s-IN�uUKPCG��ȣ,K����l���4sg�,�TÔH6|���a�|�$��?&A�����O0���t���ӯ�d�K�ڠ��B�*%�8Rp8��IW��+���'��c�e��>�����83eB�G��t�'jϫ�C�L�fZA��;�
�f 
m��}�4|��Q�Lz���;Ysց��Nf�y�sTU�b�w�����㒢B�����#���ܭ��;]f~��6a�:�'���F��TT+%�ޭ.�?EGH�{�K"&>��ªs�k�cRk{�ua��i}/ gk?(Q�e�՗��
x"�_(=̟��~3�41;A���@4&��sz!�+��Y�4Ղ9 ]�5�J��<�R0h5��vJݚ�_ϥO��B�b5<�i��sC�ߛ�r���b�=�a��&_�)8�����+���^ �;�Sb�7~(�_ �\
>Q���i� D��Ȓ<�i���X��r`��&P��TR��.�kɛF�^�2'�w�I��	���~�� ��5 KyM>���V=^�j��!��o�.��#��>"w�f����S'ݝ��J��q�ف�^�/�F�n*k����#|��ə�^{���+���~���!�O�˴������fÌ���iBX�vW�
k�W���;d͸���dV�����:ɕ2*;T,�͟Ng��t��G�B.�w	_�:�13-Z�4~�J۷�1��`&w�����(�A\jXsH��!{�(���}�j�A=���0����O{=�~(�{ZN9��{qn��B;�Ij�
K����	Lp� �o!��D��>��� ��N!M���C��ߨ�+�Q��]�p<��yB"�>��ϊ�(����5��Q�aNET�
p�Ǩ�(��>F�ܼ=7��3V&)���.$c�����R�.<CB��@e�Fkܼ���-`k C��1�T�e�q�M ��Ǿ��`��@���bTqތK���&b�>�:���nz�0�
���cx�����̌�(%M0�M*���\��7�~YWB�F[(Gu�K>v|>�S��T�񣅫�	�e�> uG5{�3zޤ�����䤅�H���b���+���g'��7���^>�'��Kb�k�OP��p�1bpb�l�h�ut�A� ���W���&l��=u-�ٙT.+����3���H�6��A�?����7j��a��O��)wH�����v���wH_�s�e�OP�!�=!1�|�T�+��R횒�y.o0�u�#<��9:
H�7�jހ+Z���e/���ũ]bd�����y��t�3�ވqR�y�5�/�)��gD���o �o��o;hy �K�=� /\��4*��<ؚ��=L�Y��=(7� O;@�\[;���@�����Y罭�r$����J�`@�0̺�K� ��9���>(�U?�!1kd8�[AJ�7WL*%X�X��hFp�~~08��}�oY��]y�u,�w�,�P�%��>��ޱW �ǸҬNI�ŠQZY@Smem6�aͦ��>��AӾB�N�8<	��ʂ�V��3��)6��׶�?#R�u�h5-h}O h�_���<^��/�����Nѓ �����=9����_*����i�Ǡ[�����k���^�q�B�z��IH�N�һ.����<��b.{0��Ye����%6;����i��6��'0m{P��L~��V��-'���߂�������I�J--|��9!qb�|`�� 7��6ٵIܽ��Ӥ_3�PB�E��cr};���B��{�w$}�M���rY�o�a#3�UE[)���䀗�t�΄R�ϱ�8'o'iě;��*v�_����+MwR��E��_(��+g�����-X�0� yr���\����{.��x*wt�����}�Ɠ��p~((�xi���ko���[�����S��4)��!�R���|������A���v���c��d�WXb#	P1�� �ԯ��vE���{fv����|K��DQgOh����y�_؁�y�R�E�VK�(�ԧ�J�1���9�w<��CEw�����D
܀V�߹���G�	��7�R�T�W��1����`"%;��2������8f����)�Wl�,V�,Z�ՇOS\���\����;1�
�����z�H֒�al� 򭐲_���H$%�ڮ�T�\���;����bK��`�� B暈��}��`�i�'e֩9#�f�с'���P�q�is�w�y{T�q��TDy�U�|MmajJ��Ѷg?�l�,��}{�w����B�}�:�j�Ԍ��!ץ6T*tʷ�Q������͝�Z�xM�.ׅ�y�~��zsHAU?�o����.g\�Z�V!�֨�p��i� v�'ײ��)���SoCu���9:��Lm=~A�uw�u�d��{��-Z�~���A�y8��¨�O��6Ew��z|у��Xll���g��F~P�oz�۲����b-�x1B��
(eޥ�;oM$�uvv��N_�/��u�	�����.uG�@n=k�ށ�����#��Ϸ���|8Y���Lv@����bgx�ǈ��.�G�.J��gEG�,��#eLz֣��k��!�K�vne��M���z�=�+�G�
hϯ�w��*�Y��9�
q���M����CM����g�W�w����2Þ���)�
Z�@�>nWo=�&����W����	, �'6�γ�f����W�9u�k?��v*�����������/k:��G��K4�JRv	k��W�oAd޾�i1惰�T��:�W��pݔ���F�����;�k<�C=�����-�N��w�Ue����c^sj&+���'i�xQ[j�l� GWZ�A�!�t�`y��K�5�-\�o O���`���@����5��t S3��/�G�In�-��.4>����[tJc������`ס
>]����/����� ߩ���o���k��ϩD�����K�OQ���K��9h8G�|!
�ݹE!���A�ݼ�/�p_㫸��|���*��-ᕺ�/�?���l���<���7@4ε���ޮ������$8	�矙��?O�����y���$��.��9����mJ�jRF�X�<K��ug��V)�[�9@��mFBM�f1���T�Yҝ�s]�^�m�:��6��6�W�#�|��&?�m��d��T��N���fU��rIu�\'dW뾆�WGvZ�g[S+� �)�I�O7^W�};��\���ڭ"K�Y����=�9�I:`��mEv�3��VͻI=I{���6�+��=J�덫�EԎ�,{��'���� m�����?���0�2��{�sA�&��{��oB�P�(ݙ�"��Vŏ=�/�D�U��������� � �b�����cf��d�fc#'��i��F[Bq/�8�-��3��w�QØ�&CǱqF��c�fOO�K}�Ț��V��<����i/o����:���#�>��+���1�xHf� fWܦ^���B�(h�;I[= ��Ag:�*�v�`^j�٪I!f�o���C-s	���[k��|j�,nP8���u}���ǋ)݂Aݗ�m�|����rv�6�G]�(�*Stv�nl_R,/%o@#L�i����A~l6w��V�����}�w�Lx]�&�;�s�A#�MWz"節?W4|��<v}q�կ=��sР���<AY�Jx1g���	h��12��pP�n�u�>$��4��pjG0���K��{�,�w�����R`f�W��A����mom�"D�'0�h>B��A�H/����^�ꀗ���
��**^�5�⼘���DwC���_�ˈ�!��7h�<�(���їV��ѽ���8\�f��JK�޷����g!���y$�-0�O��w�zǇ}@�
b׌/%Ń��8G��x`�W)Il��ՄLG�/�[`��pŁk2t]0�U�*��v�!	�U�U�@8'M=^�(�}~t�]7��_w���`a��b�@�Wz�͞áu{ �Z���h.�� �?��]���oq}f�K&��I]�m�/[ �S;ሧ+WmU�.|���������7g�b͵zR/�MVs ~3:S2���{u�u�$�o�q�t~p� �ӷ"��D�˙/�I-mqʹr���%�Kr`VՔƕ��=��j�xϋ�!;K�;,��������z���F� g�|���T��>	7�ؚA�A�������|�o�'9P���͑��������h^{��D�<mna	R�8�I�I��v��.|4[Y�ѿ�W����Rq
�Ĉ�����{���=�V/��]Y&WAuK�O����k�H���5<�v��{^���@"Ѻ�i�)�(�<���WKC_W�!߻�|��Ǆ�!?�+�hp(��N��1L��b���'/w6F��.��z�nN>�c�DߐR�sn%�`f;��8s�w�c�A\e>�wE�T���J��jSa���͘�:
c�#i�=���݅ �JV�S�l�糘���ͅ7$�_(����Xj�Z�i����@�+
���%f��	�]LJ�X��B��8s��wH�ǝ�;E
�e����թ	f��Y��"��mN��*�,1�[�ت�5`u;�!���R���oqIe+F��ry�Y˞� Hq���������֤�݃hAu�����ހu�&]�Ke�*t�9vs����ā�ͦ���1\SD67�K��;��ѕJ0�53,�5��Z6���7MV2|��&��k�q.�7�f�DAٯ5 ������E�w�[qQ��^$�k�Pׄ�l��W�.m/
�����[M�z`a�������f��Øk��wLf��1��粐&��T���ou��_��7����z�� |�""�O� 
ڰS����v63�[�!�L���-���VQ�%p}H�_��B��i�ƘA?�:����&�?�;+E%e!c0�@2J��NÝ���Wa ��������|�L.���q�%����ދ!����s������ĖnZ���F妘[�͆���tg��V�z��Ns���0���n��n��[F5��?�k{��w`�c0VyP��.ֺ���fpՊ?%}`�Br0�L1|����ݟ���[�^�Nuk���.�Ʀ0@��
zh���m}'9r��c����@��!����ͼ�>MN�X.�������e�8�n8ǭ>Z����%�f��a)�Su��H���S�:-pr�*A�'&�6�r,ÞՖ36��@��%�:K��������I$�;��ZX狂��ފ���a�!�,���k��EH7���������k�W+b���BMf��Ϭ�Xdp��~t��f�`�X�]����4=M��ᗹ�ޏ<<Tv�����z�{�x�{x3 ڗ�8�P��O�~���z����E�\nn	%�YR"��5��"�.���e��F�ma�+�����������k[e��+�2��J�ꦘ���B��4D�(��m�xЇȄ�>c�V�)���ˤJ/Y��`_�e~���t����6��ÃC��.�8�($⩙��Ӟ-�E��;m{�MW�: Mx����a�A�����a��6=��RB�'��z�ft11�_�]Eb���
����Z3!��B�B�K�ކ$(n\"5���:��x�G.Ɵ�`9+�Yi���&fh�*U"�����VF��z� M:j'���%�`���3�B��i���w䶶&P
I�J���[w�Qt���T ��^%K�T?�)��_�%�Zu��Z��X��6�h���k�&�{��Ȥ���ėX�mO��Z s�Lx���Q��ݞ|I���|�����H:���\ϟ����PhO���v�C�\6l��ᶼ�����˶�����1-��: 8�!���th�{�p�������<;�0�:E@���gǩO�-(��("%�S�q�����425~�9Qr��O� `� �֓�k�գ�y��+������g/s�{�!�ۭ\K���G�i��C���U�X�5&���������Te��|6CC�ݵuO�}�׿�|#�we+@���	�e?� ��5ݖqD�%;Xڛow���2!G�(b��)����<d��t��퓐��`�8���Q���0X~Y�� ,�Z���%��T`�e�:�������B�#�z�����>���:
�H�y���+w�)�So��E)����
sTL��͒X���}K�T7�9����_Ր��V�����X��%�8i��/�E��ں=�!q2K���b=D�۴.��a�A"CI���h3���E`�s��%��ۄ�ض�m��>)�LO�H}E?g��1x�@�	G�X�� ?�iҡ�����g���_ ��v�0���&4�Q _�+�/=�2���aR���Ue�`.Bj0��_��`W1 �5��<Q�F���O��ټ�US�/�C�n� �w@�8���ڳX#���h���PT�PRԂ�E��z#���v�gu��;�`�x��L"3 ��,xw؀:MJ��-������G送�'�욹=������u/�9]�P� 
�6�}Fz�����4Bf+���a��Ǚ�~��㞟4��4b���(+@������K0̕x�c ��ծ9���Z��1is�[ܪFi$�I=y�hEv���^��1�+�B�K6�1�v�{��>��K������C4HIӱ�ZkBjd��B�	��<.J*z�֮ϗ��@!t��^�wB� !���Ӥ�����&����p���c.�3�g ��&G�JcNb� ���񌍺ѨT^ҧ�;%J%�-y����3���v�i68�öo܃IY+��8�W9	��Ic:�K�B+�R�{����þ���Cxz��a��I�m�#�#�U��0x��n��(J��QO�u'*��!PK�a,����rm�?7�|t*-'��!h���[RZ���M�%䚸�&������p���8mW��g��e���Ez@n.<�(��2�f�]�G��t�����퍐��9�"�?�?����`
==�A�T������6��3�tq���^a2 w^�`K��h�����[�����ִo�",Y���wj0�ʤ�1�S7k�@N�PB2����w��7��!.�
K���;셉H꣼�"H��K�;�st�Ğ]��K�g�GǾ�E�D����	�� 8P"W��ٙ����	�Ϫ��_���B�a^�nl1j��-beY��t���H�	D�|`�5�.h�b��@�����}�j�x����<��"-=���(�nL!��>�V�m����i�5�tN46*~�2��.;�x�l\�l`�k�+6�X�Du��"(Xbc91gJL�?MR�V{�
pK��O��ޢ|>�ó�5��'p�C����
�xt|�����J`�T
b&��(�?U�B���f@��;�h�#���$!٫�Tٹ��3���b� \}���ʞ�ZB���'opn!��SPt]�SڬH2Y`2?i��g����/��,_�M�ֽ�������*�������$�Z��!�LQ%��'���>/��D�T��|�����q��KݤoDߋSgv�xO��u�n-<�K/4�ѱ����䃟�����s{s��!e����`a��3�W�^{3to5g 
�W�4��g���-m��"}�Z�/�x�/�S>��UC�3*0��aV��5\ɞxS�IzZX����@�1a�z}���qU�Ge��"��U]��z�n��c�B4f��n�֥��,�DNt���]U��P��]u��y�P�t�L�aq�}���a�7�|���'4�g�j�\�d[I�uY����w�!Q-�z����6L��� �+�~B�����7�Vh�M�|��&�|TJ+�٣�e��O��6���Gy��h��[JZ銂t|��j��]&�#��*MSOᤢ:��F�͏?�V7�:Y�(Ѵp ���k�g����^�������\m��×8�l��������n׵M�
�|mM���n}�����ᚧ ꘴a?)��ў+�K�5Z�K�UA���u��W;]�i��e�2�L��m�Lrp�N�ܮ5�;F��D�
r_��6���m��L���ӛt�߅�_��1���K�a�-��`�	 �q��/35zk�%�S�IଧR+^l4 ��N�9 "|�/=��� �ܬY+�/�Y+u���'��D:�o �um=:��@|}��#ff�¡8�����Dq��d�{6{��
��U���gO�"��O���Q��/�N->�^�\��͆N٢�Y�i [��%�#�={'z���V-��K� 4>پ�)���g�PѥV���ͷ���;��i��Tu��O�QO�L�]��.$�;$=��i��xӶ�u^]:�U{7P�%���8�&���L�MM����f�e�$���܎�-Ӗ����І�^�;�2X_���_ȝ�����r�h����R��x�B0�4����:�ہ���7����J����ȱ��K�0/�]�{Ig�	~#��U[���O;j����!d�I�>,ޘX��$��ל�~��B&������U����w�.�;P�ﻺu�̒_9�`q^�!q��+�W�sxB�R��h�-�F��o�6)���Y~D�� �[-Q|%�z�Ԕ7uf��0��W��U���Gw���va^�'��byeC�����s��@����V�� �=Ȩ�C����_�Ƕ>xL7��2 ��o��k#w�|�(�t�5qD�旉�0�/LSf	e���;�l��jHC���v�5T�y��@�Z����X�V�=^��~?�����x�C���g�v�F>�d�����;r���œ�T_:]v��7ӑi�7'�&��*����K��*��D3��_S@��З��͸� wiGO�yϿ���1���/J<�b��/�Y'���<�t��K-t���Ao��?��&5�Sl��qhV�,k9����������+�F�Q/�� �+;P��!X��:�k��?�_��������N�K�+R���v�
[]4k5�]��G��_C������M
�$��Z����^%Y�1�\h$�D&v�"��u�8U�����_�o8�N��,�0--��F��ϋ���*'�ޏ�Y�Y���u ��Qgf���2.��N+������fP7��yYՎ�D1�#4T񱗠��뽯�%��:4A���[�;IE��L�olQ06ya�����*_1��h�q�[oWW�O5�U�X�7��X�_�M�W��Ҁ�*�BQo2Z��ī|�TS(o2<���t�~p ��\��V�l�X&��xPk{8�E9"�؈E�#3����;Q>�k����,֙�,f�W٣� ����i�3�������Lø\���R����w�ĭ�U��[������m�ѧ"OSJ��h21M��kUop�����'C-�=#��޲�����0sv�K��+�Ĭ��A��l�6ЛԜ��B(aJ�9էg�O*J��(�N<� �Ur B?O ȁ�����-]�9`�-�%���m�lwR��^Q��e0�]�SQ�P@Wg����Z����������x�8���a�_Ո=����o��>�_ā\�^rx�J~ruQ��ƕ�ja��9F`��b��崪�C�9����_
GIT�F�ʱL�E(^e%S�$꩝ͭ�@]���Z=�Ew�c�BBɓ��,��G��i̐���T��Fl��'=?G���ۙ�5{<C�n�oM| �S7Y�x����<�;z�C�Ŭ��$5-�4��*&���P܇|r�!�ԗ� �׈����]�^f���澇�p\T���=ضK^TR�Yk�XW	��̷Y6�j�S4hr�O B>�h K3?z���7\����7��/&�By����i�b@�K���=��WXA�|k=�'՗DzeFF���L��Yy��~R�|��_ -!{9�]��K���_�8*2��]�y��_���h	����9l� ��o�Ț��ݗ������L���~+);7Ru����4}���6tZ��sԙ���|��S;�K(�9o�'���4[7A�J�����S�O��+���j24���^V�hY��|�I���*��x�:���C���m]�֍9h������t��-T�}�3�ʃ���� ��:�m���G��m_�6�o���y�����Z�2��}9�i�I��x�)�1��'���/G7���Xl0��ǯ7��_��L'W�?d��ܒ�)3L���������ӭ�DT�#�|��Cs�4�[,q�4��ȳ#@k\n2愊��, ���D�h.�rK�:�B�T�^��㐿���ً��]@6�s�#d�zǨ�l2H�Ro�Cq�)����n�D0�Z�P�f�����U�����c@�X�9��@�*���'u���R
�3��-����M��:[R���4�!fN�+��M����_��H?���rݒ�U�ɢw^�`�A`HB,g���� �*Iᢔ-o�(w�/Z	�1�'�x�:�3��v��!��5o mI����i����4�^�/W7eE�4A:x��{_���+�n)��f�3��.uViR�r,�ꁤ�Y)������V���#f`��݋<Ĭ�Fr(;:h+ ejTB¤��u�d"�p�c:�w;���Ar��hF�� ���RY�<�V��l������tx� A�Q��#�T�y�/J�;zI7e�j�V�kC�/�OE� �oq��Aq���^N�,J��Q�,'y���4z ��"�;���ֱԉ/� ����o��%ɒ���0�}>���(����{�#z��h�h��]x���!U�{�]�	�T:S������Y�̻f�Z3X�;D�<(e}�r�����_��s��E� ��,��̃^����Ǘ	���xOB��-��!�9�B���ԑ�ר����iW� 4�Xªߪ��h~,i`h�;3M>8m�2d[Q�l��BO��w�&�.�N�N�Dm)ˤR��b��>o�=�[�����b@(:!��M]$�;xx�mv���z�Mw0�������:��I˶����}���JI�
��1��{��Q8����r?���J��HU�j����A:_�'���4w��ُX�uLBIB�T�\�Ş��ϡNz������#&�
�Hԡ�̲�)�s�v[+[++QZC �����B��"�:��[�N� ��ˑrR�cyk%�D����̝����"���X�׆�ɑ2S����8��������'0U~6l�[zgȄ��X���(�����(*[�i��*��M�1�>.2�g{[�~iі�� �53`��nU�^���6F��VJ�q:�7apOKUx��,e6d���PXL*��b�z+OX�%(�x:��"��[�	����M)����/�� �V�g�8�����q�p/�c �o8�J%h�j �����o9��j��e7�Z��w��l��4��-�ݧ���;9��a;(�@)�����yMCxC����'.H�Ev��Q�J�±鄸�R����@�CjLpő��c��[�~�(K���)�4�K�1E	K{wr}-��J���S��!���E���䱍^����������3��H0���VJ���_`c�a)d�T�R��콽��x�����&e���`"/�c��:|��, 8���b��w�;$A�������*Dд�g�ኀ�G),���0�t4Z,b�*��.I[� ���mFg(��j!c55�6}� 0w�exp���cp{��;�Ձ�S-y��������|��O�|��[v��ݗ�����ٽ�\����Խp�p��Ra�m�4��x�����uc�sX���o�Iģ[=S��n-��ʊ�h�8����.�|���0��[{$�`9|_���=���ׇ��,�b�a�
��'N��\��ֻ\��VX�U;����pi�5L̴���j�3����=5� s	��e/'Ε�%X��y��m� ��l�l鬨Hu�U�{W6���8�l��۟�w����q�D��mۡ�g�_{��}��l�c�c��`������*=ʝP���ъe����Oڰמ�z��V�r�?ͯEk�>j%���ܨo6?ܚ(O�"���b�!�_;�qP�=�K��.�{lMIS����B������`�hy���j�a
85�T���v�Ϊ�rt���簐����BCk�2wG�����e���{	�-�a�1�����e����G�?���;&� k��š���]�jڍ�3L%-.W�(<ǒ�|r��ܨW����;��d@�rѫ~�M���W3B��-�կo��=��	C��F��J�kk	tȚYW|�G!%�������]�ɟ�C�\9aʠ�l�s����JTm��G�[���"
d�[:?��C��B[XyOșjDJ�M��ؖU�2�*�!����ϙ�m�|�d"1����!Q�!k2�$$Y�owL'[ ����ŧ`XP������Q�?�d���_�g@B���=�X�lF��f׵w�q�W�(=G�� !�d�J2��
}��s��!��������rM�`[�_���r�έ�L��"���n�n� ,�z�X�%�$�F�58��N1+ ���o�Evq��Ӱ�X�@�U�w5��UǍ�z*�W�C'5�[�D����}S������]�=���XWN�I��2�>'fv�̇����W�כH��A�ߕw�9��⏞�Y�����/v�%��EnT������!���(�BP��S���HҍAZ-�����d�����J��u �w=���P�[���Xu��5e��&,/�[�O>�,�SO�! ��4�]�p`x��rp#F�}�y���L��4r�Ktj����)��U�I�y��$�d��w��E�+����e���~>@��x ������a��uǱԔ��~�l��w�0����F אI�����$&+�vN����w#p���{�v;���۹����}V�L�;~��-$]���BǮ�5%|v���Ξ���]_=��?dֿD�����0tʹ/.l�/&+���}[�q�`.�J0L�G�4_��k�l��k>����;���o�$���
:�$�ǧ���k'!sa�Q�V�>$zp���d����DeomA�8�'������F���N3����̐3R�c���7|���Ɯ��wv��#���9s���A����`��Gމ���&�+`)�27ko݉h���%=�Qp][}�<�z˼���濡D�y�qy�3 W��~w7��~q0m�Z�&��L宆vqtF_<q�M)�˴ܾ{VypOx�ҭe_*���Y�Pk*d�Ȼ�C�{�����"�4ծ�b��6��s� �gΏLf�Ē��������Y?��`��馿[������1>����C�%�C�x�ӽ.�a�t*"���t�����y�A���d��Q4r���l�)X'F^q�)�\�Ǭs�LTT���ԩ�Em�ڐ���z1�o	��f;Lqm�E�.���<1`֥76= �!8��s =�bY�ڴ����g�D�,;""�6��4�����C��z�F���k�9���\�`ܛY*y�,aw�[�K%��y���u���q|�m~L$Av��*�ܧ}G�ύ"�X�>!�����W4[��xL��ub�B-����%6᮷@�����Q��G��OO���!�ę�X�l�S��.(z�9�����q��Lp�%�V=J������B��-M2y�|�k�(�1�O�e�m�2��$���A�҉X�+���b}@�f>� EKz#7�v��| rh��M��"��0�g�'{���X����l�庫t���P�㟾�4Y�����|����@��w�)�ח��vݱĠ{��4�4�lNS.���Ԧ�a�;NCs/|9���������1�Y��|z��`/��2}�����	�m��H�$�!|{���	 �lÂ˺Yt�"�&��M��qP?�gr2C&jիA)L����2$�rn�A���j�3F�G��9U�� ?Wx��P)�F�+'�p5�����?�m��h�$�K����XS��shqXe�[5�6vcҬ�r����ږM��k��~�*�@���YYq�닾 �Q��G0�&�'9��m��J���)�k�l�m��g{;���@".��5N6-�}�Oi�@v�iE�-��!�<O�4������1ˡ�-*��c���|��c,��^��!�X{S��ior�6����e��l"5��w�� �b5���p�L�f��`�O^Y_x�g�jЙ������ۋ���"��wfn����HFV}��AapeJ�a:΁��6������A�ܴ���c':�a�#��������PakȤS)j4�Ю������҆3|� K�fju��T�\��2��N�����������f�����"�OW�G�W����a���zѨ��Q�4�^�3�	��a�n��A�mm�iD�u E�!��z�|ri�r`v
�?{Xy;^����/��b�eb�O��ȹ'�w�ז��$���_9}�U�#|:>���!��� w��|n�2\�E����1��7�n��#m@"<@"ȉ8�'�/'����U ��+��������;�P��#�R�}��-(��+�����*�H����I���ݞ
5 
n�e�붯}IL&XV,3�y2�㼫�4�Z��#���#_�f>��;6�z�.�,�^+m��z��7ٌ&���0��yk�=���(�����؁gC��d���U�_�E�O @q�DӲ]��X_�� ؠ-2����#��4Ķ�"?���\bl��/��"���s����Mg�'�|��{�����:� �7l?_%�O�!}d�n�!�!!�	��4߾�,�6�E�M\g	�D5�I�1�������-�e71*%�������8R�� ?%�3T��|�Y{f�bhG"��Iۤu&������o���s����1�Yl�4^."E��WQ 	]�@UI(��Zq��K��t(�]�?��[ ������8r�+��g/�9%"Z'�϶O�~��:dZ�!�Ds=��靆��\����y��<��(�(�����fd}�b�����d�sQ/�2�j֔w���=���kn�1yt�p��)��N�\u�ABU�c�0]�CVi��U	�����ݩE����B���!MS�^ [�$�u(]_n8�����x��+��1Y�?�m�ҕ����k�z�p�5�L�c���w�����uJS1T�����D ��q��L{������ТQt]��Q�2�ɗ����4��F����料3�:�%��Rg�n%}�(�#	�u#ߍ�������j��O`�.�'� �	��RX�4��-��d��I�##�[���VSv��n�J������`�ik ��hL)kJ^�����d��=i�84��b�O��ǀv��б�P~bG����dǙ��Sg��fD��mZ�jXz��h�S�7�T��� ��ͼ�QY��WL<���V�&�²�a��t	.�e9�DѺ4�:07�j��w�q�o��l
ߐ��=����7���g��K���nW@R4ͨ��7R�ͻ�����:s�^-.K'n %�!�]3�ɣ�ߊ�q�4�3���|�~?�����R%��o�����R�����?.�(}�ڢ����m�4w����zۏH��B������5~�c�߻y d�cK6Ba_L�7^�n-l�����`{��}���1G����-r�~���Oܚ���S

��cF�X�H�E]�v�3و���#ː#y�A����@�s�ډ�JpJ��B��L5t�q��w�MK$*&��Ҋ�`�rփ��V�d����*z
���> M��&��߼�A=y�I�>�ewuL�I�Q�16��D8����Cd��r���b4�J�5�h�Ͽ�_��e��a���x� �Z�J��,�D��0��A����&z��=�պ=�kށ���:�Z�C��~!{��Ao�}���kz�q6�ٳ��88Y)I$t�I�?=7�X� �U�tz��p�
5�1�=�x|��k�k ��㓽s�L��{��E��뮸�]�iE�`@@� .""�  ŀ Y`$�₂��U�̐$QP� HΒs򯪻q��u=o��?�:5]U���>�9�ӥi�Gk�"�?�[��ց����)�]�����a�;� r�����i���"�����޴�Xl���`��m�@}�(x�%6�2�����c�����F�¤M���M?�M�Bp�	���r���� ������V���;G��-�5��l�u�J+kPڵ'X�uGFIjߎp�XZ�T�TAlf�[����1�j�&'*s #����܊d9���m82e����b�س��*� r�8�1�),��FӾ6�e,��w���1;?�-a�:{,���e�C_�[���C�/��Ye�����i�O�;�og����p�t��(,gV7�!ԭJ��s6���.�0������y�M�h�!�}��|MOt�LGbï��c���j~��1�ĳX�����z�}��Т���x�aB5��
F�;�~���S�����/�R�BL�+Ua��^W�NlѼ"B&��Z {*/�\��M�M·;�9� �v�V��q$R �K-J�o1�� ��v�۶K	���z�����Ά!�G�+ف��y�_���8�����o�����*X�|&þ��جΥ��}+�h�ZJ~!�xڄ)�-�/��:
���)�!`1{�u9�٧z!zCX[��c��V�R��x�ڰd���U�P����&���ry�᎝�@�A�"��hf���9��.���Y/���`����$�Juگ�/a�d ٻ�w^t�	�|��&vH�S��A�޻AldE��_���q�0|��|߻n@���M�ⵯ�xJ��⁂���r�o�X�)H���F>���8hMt&�ӿ���ۡC�V*��m_�[�d�K�R���6�;/���Z���י�Cl�����FS)�ZB#'�\�ָ�f׏��1� �w<k�=��q�(�"e��|�X>�	����O���D�T���툴�.���D�������2�j#�@��o��!B��z��N�ހ�˥�,A�)@4����s�/�X��*ܹ£K�p�b�R�,����TJV0'�x�Hk�ol�w�qY��
`%�)�";��e��\�ǌaK�
�׼G��/Q{��L)g�.�u��~.��o���#������&�iTZ'=�=�x$��$�v�m�(ǰ� FM��s`|��q2�A��m�M����HM���bam�dk��|��[�%v[ß���Q����o%�컗�,M��c�;(�l�M�MG�d̪O�;�ZQ�G7m-�l���K�c��)�>k�Z�����)w@>�����=�	��{`ѭ�&è�Kzo]�k��|-�e%\g}��}̡Je�^R,�M��,R_�=&�r���ĝ�����/�"��Q�U�6c�4x�©�팿A�����C���A��M����+�x%��6ੲ�hn�F\��y�O��b?g��N�a>ݲ�{E���~|�������CL�&�4(-H�l��_�M[Y86p�����:�Jb�5�a�p�-}m�nL�{0�v9���_�jf���6���-R>9b���>w��O3�O���@#��,��3e#L����l���ZP 8ht��QȈ�I�7@����ҕ�A~�A��J����,���Kej���PJhilk�����Wt]~L�l@�1��e/����b@j�J�L�N��8���S�)�Xk ~�� 
�W����cX�tyG�������dR����)x�œ���V�<��&�E+�M�@������S��Д�m�ࠆ#f����\���C��7U ��2XJX2�1�]�섽�<�X��XJ�������H�ϥ�pཱྀ�O��уR^Kԁ*?�<������ �xi��!�q����������&���/5).�x�O9c��~�]&0]��J�o�#�����{Fd��J��Oc'�@D�j� �F��{<�.ƙ�X���E8QE��T^j����m[��,�ZQ L+�UK��A�X�>˒E�Ya�Z�ne��
aw��%��YI��2�CT���\�Or!s�����ۍ�@�{l+'��\����,zC:��z&q��?R�қ������(/���XTfZ�N|����%�xU	(u��-h?/;��� ��c2�!rM��~����Lx����3�=��������6���ͦP�� ��(�]��jbܙ�݆0̧(�E�&��[�*���y�����aK#'(h'z\�73�0cs��G`0t��Y:��S��~CL$,��RȔ�^����G&��z�Ԕ'nVZ2��niT��U�v��&��*� �#O=!�o����c������׎
� M�e/T�tI�n�N=��:�~�Y'�����}��c'���(O5Y�;��D"kk�����S9[q�
?3Z�H����7j�b��}�e�7��#S�R���K�7����և�g�C��r��
 ���������`W��9��Pҁ���bsk¹��-�lRx�cv��#��L�����OY��æ/����l:Qmz뚓��B�o]j��U�6+zq��|��W�<0<��m��$�3R����	��쐢��?���ڷB��j��9 ?� �!"]Ʌ�Cn��p��%��e�KBAs��cD����nc���� ̐�	;��ݝ�j�H�Ch��@%���J�l� &�H�ܴ����i�gj!r���J�
Z��2s�[�N-B)����|�e�N.�w_	�%�+Ͽ`q�I�Z�e��_`�J���D�^}���ȯ��nkPY�nV��m�d>V��n�n36�����N.�=@M�����ޘFl:�&�BX
p^�>"ŠN����	���L�^�R�Y��<@^��H���oT����6K|�=�xʹ��l	F:�1~���",�G�g+��ȝ�0��=�����k#�U�T'��^��s:Ժ���U�� �N�T#ʚ{9��&RC�������Î�Y ���[#z�Zb6���[�5�����co���w�6<�`���uE�i���`RL��	���}�%�ݺ���� ����ODB�;��[��ͪ�����Kh�h�ws!�t�ZK�_�p��4GՓ�b&�&$�L1�rB]��T��f�{a}R	Y��6�n��1��A��gw�y�A��?!Ƽ~Z?�c�Ύ$�Uկ�����(@E��YAE��,�j>�[���g��KQ�%#�Q��_�a�I|~R4�0#�M�~?�F�.w�.�?�F9yU�A�y�%Vxze�+oY8/�y* ��n��G��;v�܍A����X���L�漜:T(4"�k��o�\���$w�~��2�}��|�M=���| �u��Μ�Y&y��VD�&��W�����O*c=y����{��Q���$��:ӐM,��8��k�m��h/e|���n�K�*b8e����-:L_qAE�5�4,��j��K�7�N�Q���m���H{��P�M���?�v"}��f*�Hl�Mϥ)����P�P��3�7�pB��:�,�#�E^g+6[jϸ�}���]�|v������/؟�<�T�����uK�x:&>�٣��YLP��R���eS�Y�`���A�X��L�jn����4�r�!\B����A�Z�m��,G}�k#�4c�f�i>�E#��W,3O	�Su����I��o��@�i���z.�uO�r�C�QG���0c��9🭒.\�����5�UG���ɨ1Gޗ<u�g4�@K]��<Z,-�eW��/�-���ǫI$��c��J�<�6�O0�nzq��_����T�U��ѓ9�Մ�n�O{�e���}�A�����Zb����ǡ����H�n�p�v7�=�~�ȧ�ϴp�%ԭd�z8x�E<w���_CJ��Õ�W]|͞�}�l��������>!�n�Jw�L3��n�]C�gʍe�W�,$��C8q��x�`=��ĔB~��(lX�2�����}������>�߇�������}������߇w��&Rnh͔n�_��IV�{��Kg��b���O��U�wM�7fM��ow\�tڞN�(1��V�r��Jz<Z�����k��+��k0��a,�A4k]��&G�� Nk�>{t�C�V:�gyA3�#}ETv����f����ؽV�}o���^J�RS=4����[̽�7�3>veJp�S�TM�t�.8[����f�A�2I�q�н�IU�2�+7W��%�ɌoVʳ,��//t^I��6�6?�>#������4���6�ʧ���?�V����L���cr�-�}iO/]�L��ط�����<|=j���S��RB�=V�`�����9wbO)���a����o��������$��G�0�J��O���g�v��y������ �, ��\;$�C\"U���rj�	�,N�?`'�5f3,��.şX������R�7���^�;�Bh[�{�S�ŏ�p����y�^���zU���_��8[��~�m�m���Z.b��cǿjpGr'Iڼ��h���0X.7�Z}��fn����ޝ4�J\|j�"�#*az�+9�\Ò�y��vM�&�ZW�j�l_,p	�Noۦ��oyf;���t�Һ����N�^��0��_bʵ������il�>Z\t�'���h��ө.�tO�z%�H�
p�d.�B�z]K��#Yo�ɩr�h�ҎBKJd
�Q���e�,M��=�[�3,���F��ќ�g����"�x0��위_��^�O+�7oڌY;A�^��F%#wv��.�`�ǹ|�7��v� 1�Gu5͚�Ф�}��2K�J����"u�PO���#�Lv ;�"S0n<a�Ԗ���Xӹ{��P�d]���kp�MaW��,�Ľ�����u��[(��Mر�7D�I>K_�y&/���c�j�q+�OF���Iuqj^��A_��5�lXa�CZ�dh[݂n�	�`�5�$��L=���H��/-22�K����+Nݶx����8_�5�.r��=��nh�_1�6~�N���w�P3��*�?��p�2�8�a�#wMU���m�L��p*�mwﬠ0�0[��yib��a�j���4��8��L��v4�4�^���X��m5=�$t��13�^�~�o07��7�k�}���y��]���l�,Z�u&�o6�&ee����>ʒՊ��V����r.�Cm��_g�{%F�g���32l��u[���'������C���j\���%��X���3lZ/�n^�uIzhV#�\����*Bcm;�4ܸ��Z_|6���,�|�䎷�)��`"נoIQ�b��6ȿU�1�C�ں���~'��BЯ; ƙ���[��9�%�a���ř1�L���_���}i���18v�_�e�\-Y*_<�;���oj��a���r��ݕ^�e�M���I��n��q�:�#l�>,5�W Y8��挡Q�9�>��_����u�Ƹܻ����q���sM�$�2|�.����Q���w�bNR��7�Du�Ǽ��z?Z�l�(ꕵ2���lޔ!<���R�H@l�)WW{��	|m��y��FZA�dn�K��pi�<h
3>��v�������+ղ�}ߡ�T����c�ϑ�֐S(nmVHjN)ƫ����b��m��vJT2+� /��&�k�8��7)S��[�\�a���4�[�����lm]l��6�<�zr�X�x����x�m��Ya��Y���QMN7�V��s�t gmHM�@�xJz4��m��G#4�����HC��FG����ik_=z��������낦[<�uZ;WÉ�&�96��H�TZ�t2�j�m�)�� �����}�#�"�����^?�=�̍�ʍ��[�qi�8o�r�·�P��w9�	k���Ԍ �Ѹ4|]`k�lu��ۋ����%f��YSL�y��;ȑn�q9}=������1��}��� �Uk���q��-���)��<;�����/6�'�����h�gId�۝,�_����Tb}��&�]^uC&�4�����©Ǒ&7�c�����9��V1��חT�tN���c� >�й��&?ߨZ��)���G�nd�,�����'���/z��Rh~��R��M��������o���	�նj�qF�MRՑ���Z��vi2�Wejx�*������ :�{���=E��[�ήܚ��'}�D���Ԙ6;�L33̽��1Wh�څ�ݶ|���\�`^n����!e{h�Z@"�'!B��H�B�C�0����I�cT׌cъx�{l�k�
R�<��sP� pj�w|ݧo��$=�_TTy��c06�.k�%��G�Ͳ����\?�H��,:|���9[59��/�5�w7����)oSeL�פ޸fK�c�6wߟ l�a�j��V����?�a�p�9��Sd���R��׌R� �j3�0�ܙ�/i:�L�� /�l�X�:�h�ɇG��9������t�믿�Z�L��-��c�[U��}�<1�G�<����\-ێ= �-�s��QI�a2d](G����7����N���M�rJ�g��� J�ހ��4#n4d�H)�m�q�����A�D<�s! HB��L_�hӉ&!~z&�TԍE�lq^󣒓��΍74%;R�Ǡ�k6t��gMέ��k?��a�� �R��SMVX�ä�د��f�!��b��B�֑��Iʛ4�xf��)��������[᫦%��[���H�@5��S9x"���x�uk��7�D;ܼ�S�u�����$�&���������j!�.�@q�(�Mp	m1=� �A�m��W��^0�W�m��&�1m<�;�+��/��˄�] �;�������H��4ܑ���y`wN�/J��yyf~�[/(2U�Q���~��[j��ЉOx�l�ι�ݷgj���/�(�I~)tnq��w��y�Rf,���İ`���5���ݘ��uN�"�Ó�u�L��L��r�w;&G]��5}�Ѝ��Hl�0l�O���_,���H�T�r��S�7A���͏W��ރ�V˝�_fb�uhx�!���*,���D�Fɘ̤���X�9Ob�O�fY�y_��?/�h}3�*�r�=�8��J��^�_ev��͘���y�u��?���v�@O�|�p��Ə�\M������:�m�-�W7I�6��`l\T�n�:�4�rWx���P�Xl;*�Ĭ(�����=�����LlK+������� j��ݩ��7�-]}@��h����+gx�2JڍS�P��4��:o�ju�oB��d�aoF�N�n��V���ߦ�>�l�=�^�W���3'�>�40�����K�U<��m�ٱL�s� �wӲ�WI�r�/,��ıT�[TA��5g9!�)v˳i����R��N�6p_ �'N�դ��x����ϔ��M��
se�]�^d�y�	�	��e����m��c�yw�����A#k�7IJ`��/�����k��^U���9)սyST�Y7��.��J�s"�.N���� Z�ĭl��"��&�A�^��ç�9����盜wv���ݚt� P6-M�s9�������r3���_���������m&ҙV�w�.����B��m����٧WV+m���M��!ϭ2\q��@�v�1�Ⴎ
�43s�O=��|Y�[�������+�g{��\Y�����
�v�+� >�8r@V5'�a@*��.��s�ƚz�����dZ��j�Tz���/�4��L�����(6���x	��5���Y��2�=����r������±�'�w�W�� y�ܼϻP&{�Z���l�U����� ~�EB�˩����fh8�+a+(��Q.����VJ���C����_I#��4�}?	����,A��ͅ��,=��ձ�t��2��Ykt�zCɶ�P�:��6�Y�9��`�jz��/f��Y�nFX��J�	��Ǔy�λ@(��$ ��)�����m���"�?PrKٷ�;||��9��-.��^��&B��$����s%�����'��V�ra���� �R�$�q�M�:�,:��;�b9�\K��i1R�������Qg�	a�Rj�ə\�K8[��o���n �X��ej|NCQ^N]Oy�Rx�[����7%���P����+)!�?�0�{GWI���$������e�eZ#��#���9��^��ƴ.q�1'����^�h��m���]����z?n��ޝ��-Ե����>S���)�m{�ȝ1}����	�,b������-Ԗ���c��__�ʘg5���Lf8\a9��6N���k_q�CzI��8�I���""�`pj�\+D_o�����������E̸2?�[���D��fC
��b*��+�<X .�\�5P�:���O�S���oj�T�r=0U��>�+���0�nEi#݆��h�_й��=����;9�)�QS9gr-�|.���u�ѳ�j݋��tu5t�i|��ƮhI%�I*L�s�s��g�9yb)`ƣ�����GA���r�A�`Ͳ���{��Z't����p���/�	_�6֧Yav$1�@�:��-�V�8v�M�1Չ��(P qn�]�?݀^{����1K	*h��`�����$�
���yS{�^��u�T!�5�S��UK��:��[R���ή~ �dL_)j���{�Bi��[q���?�8����R���?ٕ�CKb斃?똈�,iđ����s�)������k�l�a��=��"nN,]�eZ~#��C�!��F��p�1@#�M�r�����I���������BRϮ�j{DBE����e_���e����h�u2�P���Q��
��=��G�d����{5��!ݲ#���YݒR�Қ_�/�b_���?��#��&���
��RSWcb���F�G�����L����.[e�n\�/Y7�Z�?���=w-�u��~��RB���R��G�5�z�HW׬�:�ʥ'1���Iᖫ ��Mɏ���g��=!�Bl���~��OӍ�H�Փ��>�=�q	��ܿޘl�'�C2�֢d?�N�p�Ǔ�����4m�οhu����~�
j0�,F�)����'gt]A�<�B6��\eU�6�1v @�~�����v�:	�ϝ{��!\";��'p�ΥQ:kA�[�{��ʈD��������x`Zݛ�Ni!�-��50�Gx���N�y���_+����%�o[$3���P�����0��h��8�c�����f� ݖ8�74���`{��g�Ǉ��Z����6��g��C��Ԕ�ICkPx)iȬ���y����axK�d�	��{�M}1 ��Ĕ�\M�#s�_?�~ez��s��C,q�j���K�2�prR\�k��̹"|9��NZ@�PO�����!�?��:��?���ӂ5
i�HZ�{���c<j�Fx�WA���1�]�9��D�ˠ��jo+�u�^�������O�v�aZ�����P&�zAZ��l%=	���x =�Q_m�ǔ]%��ߖߦ�c<��Ah)��-7��M�>^�#�?���+E�W+��Y.�R�5����s�T��UyDUI��T�t5n��0)T]��
E����Q
�o�p���/S����� 1:�Y�\_#A��2��[�%�;K��@�p�����r��#TV?��!��������@J�q���?2'�U��:�L�J
N���a}�b�Jcc"B^�Q�/ܐF���+cި����{x<�XL�V��#!�I\�������0s����=����a�٢P����Ǐ`[�CO���,���FY�(�y��ۛk	�1F�ɑO�N����#Jv����+�3��m%s��#R��<�⚋9K����������U��ofq���߉?LK*���K�ϑxQ���D�h��L���ui��]�#-"��d^�e�~�D��۾I��b%�G��.�+8�ߪ�Ƌ�3bq��<܁�\�0imw�!"I�ÄI�0�u��.A����u���C�� ��Q�?8Q����$Bw��:p=K?�iW]@��mq�B��A����F3s}et-G�ú`T�g�l5��j@�tw�M��
�J?�yh��Y�rGF�:�]@pGC��Zo�,��0�,��a@b|�p8RwR��aT�W~o�>>��@�ړ����uS��J~��M8&w��+~��?�p�;�t�h,lT���t Ը*BOR����;�C�AY�����ʘ�X�[�nX��p�@2Zm��W�S�3�ͷM�. �Ø���	�s.��)��CZ)i�9���5�f�D���F"��c����ŋ��~.�Hs��2b�b�!͑�����l8�`=��+����*`^�#��o�.tz�����m�Lm<{-a����J�iKL���%���'�/�g�=jP�"��1��(�Y�lm8�E�罀�ĳ `"��tR�٦�{�b�It�\B�]m��߿[�q?�ǲܲ��z�W.�� ��,�\ind�%"��W(zAC�B���܎m�����¢�;H����V�h�������Ѷ}��'���c���m�&Ps�����Z��Ыj$o��Jb.��N˖a��zp':������ˋٞD��7���3b斜�+1��Æ6�0q�V/Ag�L-]ꔇ��^Hc�}u��mi�v�u?� ɕ0�nȻ0�(
^��*�m4Y��BPY2��bDЎH,B���RJ�5&�X�Nb:!�{_�|@�'�@Q����B
��Lb���Y)=�;Ψ����@��y��b���Ao��f�{��ό��	�k� �k��g����)j�YCƇ�h�'t���ɫ��\P�䤅�Z�精	�'s��$�&TF�Y��R؅����`*=��Z7<	?�ڟX��N�����.����G��%�7"��ǐCV�X��M�ʠ��(o��F����[ �3�#��t�7%�b� ���zAm])�;�;p�"eK�9�E�| �� [������K��>����ɟj:��5�X< ���F��r���b�ϕ)�A��0�q��J�&�#��
?L��Ϯ�㳮gl�|[t��2�������ϦY�ƛ�L�Bn�dV8�0�X�'�	w���V��F��a?u����K��	&�?;���!T�� &�CD	�겆�Oi��0�۲�D�� +W!�ҋ��v�D^��}W9�FRl�!����W��[VLv`lII�2�,^�V=�yJ�k�g2V���L��woF� .��+�ͪ�a���}v>�H�^�����=��?ƛSeB��w���GMZx~| �{�����D/��{�h��v�\�_�2'�{Т��oXu��j0��a� �#k-x����7��Q*�����(o�C,&%���n^H���,˄���>7�=1�;��$�J� )!����O\�G�C�xo�ƱcJ$�<uC�����VB�k�����S;�@�@����In�v9訟�<)�9}�޲r�g)�kG$�şX�;�j\\�6K����d|��я�'�8�4�peO�S��ߢ&q���I��O�G\ѝ���}�l��_p/��H�O��/�Z4��(�x�tn��`�'{<�/7��W�e�t�*4t"�D�����<�01:!��G
R�z>��ȼ�\x�h!�a
��u�K}�d���ƚ.����ܡ�}aK$$��~���L!��L�?��=V��x`���D��:,�+1�+D�Ê����I�<;��caN������(��7�Ԛ*��F���.�R@����D��,J\��2N�^$b��e�s��ɚ��K�ͽ8�;�p>Կ�ၩ��( �f���sm�+2WB���WC��W�4��)J�&�� �ڋu��.�c7�����0R��:�|d�L2������ �wm��}��E
7ܙ�#������������!�O��e,��b����CK��yc�`*b2�!z{�����@�6���/��m0��A����՗�y��Z^��Ⲣ��ϝ�\n�<r�)2q��^��)�a�5�V T�ܜ6�)�C�(��Mb!lw!?U�r	8?k�#��	�=����>��r��kU����Q�Z�g{Բ��[�x�]v=:�bD��ҹU<�����7���c�rɕ`��{ȜY�B�ܰ`N�_pHCs��&a�X���ER�0��i�P��A�sH� :m砵M��$2��W{�1�j�nz�?������������P;��ϪJ$���;����W`��Ӣ���Q���0���RƩ�R�$�\k&�;dr� �%�=l\+����&X�.$�F"P�s�*D)��}1����&�r��˩�9������	�����b�D�b���4�c-5"H���_�M�q�&
��k��7	�����~��Ab ޏ|> �)j�0�����C@r|��D�^'�;P(b� ��?ݾpۂ.��t�zn�:�rd����R��dH��Ȯ8ul����������5�j��>�?m���N�_B�ٽ}���!ma��OE%
M7��j7!�]J�m�t0P�[�%��T� BG_��Z�M�+�I�D���F��&��ԼcZ䛸(�1J"_&F<��,��r�N�O�Kao��-Ý4���?��5|�<B���a��xS�g�����9��/M[���f��U�mڌXn��GY���׈���k����L�/�~k�(���w	r�Dδ�4P�U9���	����i��Uo��T�������#��b�����<��&�`�Fѯ�]����-|��q6��J�Ԍd*&Z���"�r
'����$���ɦ�σ0D���d�GM���"d�_�`�-��%�a�*7%�\n�iɔLW��� g��AL$a����294٫���%;?x�Ʉ^b��X�}��@��d;~WW#/	Ӱ�JV�;�r�3�J����Y�`n�
�$��
�DX�'~,��É��>�ҤK��%�e��A<_���.	X�@�q��
��#����k���`�qph^j1䦠������绸#5�x,a����)����{�[�qj��C�߫�d�����\ż0
���Ejv'���b�Ȍ�*�����x��L=|�[�8xD�=B���׍�c.sq��xG����e�]X˔��_�����2�@�sd��%���Ǽ� .�3O?�/��J�ﭪ�,�ݦ[�~��+5����8�b�U
�E=�$j'c�h@�B`-|+�r�kq�[l��#ۿ<�_������"���ͪ�ck�XӇ�6�G�^at�;���OT���,��KO�������Y�I{x�/B�R@~b�K82�W!gL�/I�ו:%�IO;�Ȯjg���/�70�^(�ͩ
{���z�7Ӽ/߫��m/�_�92�i���cý���m��V���q�k�&Վq��Z!�R�ڗ��[)o_g�����ez�ԛb�]��+��v�s)swv�5��q�d�ZY��P�ԭ��6,�
���z!;"��sl�⑌:������,V.h���s��->�V\�뭹�8͸	�����♅kӵ��)�Z{�##�&sii���p���X�n��X��5�pA��M��0>i��ʬ�d1�e�s,���\V��g��[��U�l-���/�4��FgLS4ѵ�QU���Kvd���EڬI��g(���.ɏ��J\���p��Y�tlؼ�џ���:������\]��CMuVj�[���g8D���bV�#0��o�#���v�Am߿��B��i�����J� ԬLp�%�!�955_� ��״��_���ްG��l�>�w���f?a�S�ݔ��䛌����ڂr����K6_�/�eC�������;\�'�FV4ί`X�.�&�H�	l|Р��}�R !rY��[������P�ȧPk���*�����S�Ғp7=�9�{���ˍ�yOf�zFSs�{�i�LFG�\眇���S�	[gQ���¤\w"����3�Tǎ�[�	/���H�G��|j��P�|��?KI'�z)f�5�(~4�����{f~[D+;�Q?���)���YD����&3e����y�C��%eU�9�q=2Y��O�iM�f�y�5���̠���nB��/0́�܋q�pR���t+7R�EAgO-v���}m�Bg�|7 �"���GRhe���C��lv]�90B#Pf�@��v�+3��`�ߐ��B���������!�C�\7Oa��Xz�{���O�+UУ9x�|N���	��V����l�os{�WŎ�}�
U�;R�lN�Tu6�ǛBw���$8�X�	�SL(�a��="}	ڽy�Be�E`G����4�ФɨT˥����-cm~���X~~qR�ͻmOqu�R�S�/�Ew2Tʉ����8{�Lt��i�w{X\֍�(�:Ư�/i�Մ�/�MlF�E.�5�F�0�h�/����;����*����MvRc�c�N�OU�� ����n���)�Z_j�q�2�jͪ��TKd]�e����tJs�i�_I9/:"a=]�M0�G`��{�'����^����O�>V���
��(c,1]-'b��s�W,�d���_���a2�q�>�^s������
7X+����&�5�:��eW�B��_�J{�˶9���4.8��-�g
G3��d�y��;�Uz�:~�n�]},�G?�<���H�f�����,M_s��U���>u[B&�������=���i;��k��6]u���)�ջ�l�X5�ݹ�pu誱�b�;l�y��gD��<t���?x<����꺧1���>A� �5�4#�V�ط,��.��xE��XFM[ް޽Ŧ��y��C�����k�u�eLs�һ��r
���x'���^��fq~p�f���Ma�X�:��:���KhNmb������=�}tsݡn�
����ߏK�7}���ԇ��?���A~��|e�����C7X�ikWl��������hW�������{�Aj�m��zx^7tnR,~��a����Z��N38j6)�;�56p�S�,+7��b�ji���wy8��9~9��n�w[��D��id����O�)�n��jޗh����4i\XO� �������&�
�Y�����x�Y��8Aw�u���a��NPW�L1�n���8�Vڧ����>�D
��3/�^0�
9q�x�\���]����9���`�)�29K\զ#q�>.ne٨Ñ�7���I�Vs!j��z�v]~����A�p�XU~��� b|�Aih�g�ӌ��{m64�s�5/���,�����]��b�{;�6��{5=q^rQ��K_�-�3#�^�/�Z��PM!�/U?�u��"Ͻ�'�n�2��r<�e�R?Ԝ9b'k
��ճ�м�m�Ӣ�G�[�H[��bw0z��n���)v�M֫EۧT�&�7\�ʞ:T0�v���rs��u�%��|�2=4��y���3[i���t��;ÉO�k^�N�9N��S��R�|��5&������͋4	��d�R!Sv���������g���mz�o�gʐ�MbӴdSD�?�_����A�:��ڝS��3�����8�<�A��Ow���D��*�����p����;�Yy��<U{�~�c�d�!��9��cҽ�d�)=F��!-c�{;/�ջ:���49��� T�[o���eSÅ�zǙ�a� �U�ѱF\��I �4ިZ(}�"Llz/�Ȓ"[��н��S�TvM�g���wS�:��B*�w�.=�d���$JK�~+!��� 0�+�m����7�/h�G��u�������e������N)΢��A5(�E��Ŋ�L^��h<��I;�x`םG��;��f�|R�	�pbo8ߝ}���l��m�URvq���gw��8zr���hR��}?q����{�e��p~��i��	p�eS*g��?o*�u(S�n*��Z�Ul�m��^Hi�񸑮Ա�[S����u�w�NW8�;��'��=r��W�a���;4�s-�t�ݸ磎�o�LÉ�� ��1ç�m�~��Ҹ���
Y*ˣ4�������_�����!���n�������ğ)߮>�+�5���OD����l���'��}p������N��I���)�����.��+�,�Ub�ZF��VW$��i.��X;�~�Szm�U����.�>]�i�o��ѡ�y����G��T���[+��i�'z��a�����<�!G(x��Ū�xG�k��*^X�&@_�$��Pt�0��8�{5�sR�ǟ$"ծC׸�(�53ڃ�B�^U�׸թ]~�r�G$i�)�'$A�z��e[��@��t�z��/Q�������v����h/�K�ߤm��ҀMX��瀾�?�N[9[K��/P�o�n�R�7��[��]� �-��K��cqzA�G}q"89�UG	�u�sTuu�wX�Ast'��h-0�o�Qs�5���4t/���-���r0zƖ/���ǲ��t׍��	c�FZ|�#;a+�Q���I�!p50��e���hX*ҡ�s�Xϛ�^��d����|=k��B̶I�;��ǥCِ�5C�����>ơ\�BԸˌY�:%�<_T�EF�h�x�&�94��J���Ɖw��u�<Z_�V�;��ķ�;�9�ʍ-Z���0�'���< 4�
��Ӝl~���_`�>M5�ۊΉD<�V}?��:~Ţ��i���J���(4F���a����5�VZ������V�i}h/���R(�yz������vd?��Y�����t��jRS�N��]DX��4��n�~����=O�*���C[��$�"����}R�d���) lK����(?waZ��4nͩ��K���������-���P2����:fC�(�\Q<d��~Ul�&܏x M��;o��A�AL��z�(ԱO;¨$�@d9��P>l�w��e�ａ:(���%v�'սD�OF���&���F�`�\:ۛZ������ۚAu٢W�����Z��b��n)�&�4q5:G>l�!1�e>>3�@L�M��q�@kq�@NU�9��q�
ݻ��T�΢�>Q� ,� D��	��k n�Ũ�àob# R?%-��[N�'��Ҥ���!�*�u��߃�Hz�1ʕ���r�2�{�|��l/���o,}�|�5ѪΙ�hz���g����ub1(��8v�#P�k�i�ʐ��{�xa� (�k���v�B��Jb.�����Ո*G�q幧C�x��n�&���=w:���kW�b��%�E��ɴ{Y�����K!�����cHg^�J<�yo�o���nY��+��
�$�'W�����£�� �?I�싶T�!AX=G�ۈ7mN������t�!9�6�"D6|�A˔��H "�(0܋�7~-Q�Vʿ&�����%�RV��J��5U���{�Q�m\��$�E�;��*����T�*��C�",����q����-w�Q�Q{2.[=��J�a�y$��v���)q�~�:S�T6u,�T���{�����+��2�W��D�`$�>ܹ��`�7?�����y�K.5��ࠔh���˵��,������_IW/Z���(��Me2��<�������Уڤ4E|A�eU*SQUi9�`��s��i�6qT����r}��̫�(�(B�~�܋�}��ԟxl$�8<o����}ښ��#7�73�n�/�ә%�H�}�МG��2T=� 26MQ63�[I8���ё4M�Q#-��D����L����*3��݄z�$m�v�W��v�mBS�FZ����>I����U\�j��Í�$}33CC\�1���H��������|��7���ER�m�y2�����Q2��� Eb�K(jE��hW�S�@�� >;~1����ĩJ��fd#��NG��� �x%��>D JF"�4���p��|��*�՟���A�p1m�I�J�r��pU��D�B�����?����m0ɹ���Ę!;��~G��k�v���8��1wFm :���f���!�����Q�T�I��U�H���{.��֦nk'��.0m��#�AO����y�0��С��}�gq�Y���vj�v����,��.!���+��E�r2�*�7y�F�ă�*{���G�����kZ��چ��7�9k��k`�>�]��K�
�s/���K��wA�/sX�6��>���(z�8�~]9g}�Q[#�$���oюNb���+�N9�0��Qf���������?�ӄtézu���-o3�Bn�3T�`̽�te�������=���\�&I�
G{����W�/��R״6�tV��O��O-�r#FU'4���*?O�5!�Ώ7�Y�(����pS��'z��̏�k1�p�ɑ�K�o���I3�������� 
gf��$<Wr��M�����49�$��	)�����~It�2��3�{�)�vB7@�7s��c��a}�j�}�ct}��4m�VgV4�C���_=M���qͿ0�L�=e�V�YN�ϫ¤%��`[F�A�0�g5}Vg�D�W�����,]���ųg�ߖ���}��gND����%}�3��"<�e�b80LUƮ��HsێȒ0A��B�0�@����Piᮻ�N�:zj���u� �� ��<f)��I���n�þa�r��0Q�6��%F+��o���ى���.��h:����?��e0��o�OjV�e��5��ǜ��)W��)~��LM�S�F>B`��������pj|���TE'�<I�%8�F����-.ŁrhtM�bD�k�Ku���2nV��u�� ''Ck'�j�z���,��"����EB�u���{t����,���,�5��cN;X���÷ӟ^6VU7���!���d��CX��c���?�����=���6	ak�x!.����-
����0M�9o8�#��"[c]�K
9�.C	[UV\��e��"x!W�:TF������l�9*/���D�$�4�*��BDmP��	ߠ#��S��N�;$��4nĨ��A7DIi���ش����G]'��-�B��a�m���K1� Lb�bB�xz�~�8R4K]��=�3ť�Y/*�0M�Q��'F�{c\o�zbِρ�qU�s\�Pw 6\6���ھEou���(�wbZ],ձ�SN��F�hY�f����sy��e#>E���y<���k��z^D�~]F��e4�Q���V���<�y
6�����k�V�l\(u<ޮ||�Ky|=FLڏ����1�GKk�q65П#�,?~G�Ԩ�#�Qb�P�)
ŹzJ�� C��Z��{�k���;��H�8�6�񾧉7w�  %� J�p(ŶV`��p|e(��8J�������y�X�k�������֛滜�܄�v]Bu�VEU���dЃ�	﾿I���@�i|� o��燲��5ӈ�J]Jי`��F�0���?�K�B��R�4E�� ��1��k҂���0R�b�2c�-��|:�.�g~*�Hs��S�N3F�V�|IF���%�D�F?�ix�4��ye>�X�8��&�(6�}l0��>mǂ��k��2��܌v���jdx�=F��������D�֯*�5��d�}<��8;���oG�����=z�
���6��?4&J|����a�!Xȿ�� )�6q�9�{S��u�Y/?3��E�/�q��ɭ�tt�����&��W�E����
�".�e�E�( I@T�����H�*A@�� 9JΌ�䠒��$�9����n���Ͻ�TW���SUӓq�+�0����@���Ը��o���෷-�|��-���vO���>�԰�T�%:��q
�q^AQ�=c�m�}�]s���7�#w_���	y~����
ާ^�q�B����x��]�@\�9L�03+�*��n�����Zh�uw��;��N5�f�J���'�9�]�|�Q���rT�ɦ5+���wY�^ �U�߿=J�k��rW����͝���K��v.��t_8�s&��u������P�.D�8�t����{�����OS�^���y��_���S��}��7����?�^9z5^�E���Dة�|׍�.Y˛�W
��++�.:��2��A�د�ةg��lվ�n2�H稍��&	Ҧ}�3�vg�u(m}�@�����Ř��N`���Fc������n�/�ݨ�A��,��z
STb�m~���ዛ��r�7k^�v'H]��ɂ7кn0ts�E���5�Ǖ�qu�Kۑ������,��l�Vwk򡬂6��4ӯ�o4B|�j��'�#��v�g�'�v�v�ۊ�)U�%"Dc%�d?���~�Fu�!Z'���Y�i��������}�+���%����ŝ��s�z���ʎ�����3fu�y3ЋjR�p��>�PM��mZ|�Ӓ~�G4��s��/}�XB\9��?�\�9��!�hy��gk��/p؇d_��]_��)�ZB�&���#Z�\�dZD�iKύ ���}0���T�E���Mk;D��D�_nw�������s��mY2�/<o<h��� �c0e<��h�M�FJ$�n}��h1�����(/x�i��!Fi�:�����l]%pcPDO�m�H���WH
��?X�.�����_�ig�����}kR�[�
�� /��y8��E��l��4+��w�M;�x#�f(wluaa�J�.�dbxn��4�����2z${%���������8q�����d�*����O�5���n�;�O_|�{|L(�X/��`(��b�ͪ��j{�T�L�'�1S��EE��Y�y���l7Jn�	��˭�k���OA�t(�>V�/SCS׈4�����q�7��,��B��6���I�Ш4�=���.+�T3��ZE�C��?Y6)t'FAL����uDf���W��R��=�S���M����tf �S�ЎsRV�SVR���C��A蒇M�%h�S�ZO|Q��í�e���'����@��p�ֱj���cb��ַ˭ϟl��2����h֗�;#-R��#���P���� H�e��1��ц����׭5�ow��	ʏ>w��u5�� �ho/9���ZJh35^�܏���+�)7]}���;��o����:��)h�M�c��d��h�Gtv�[��vT:��&�5�/��0�^td1{���N�f��)Q>��ҜMn����ֺJ�h�����8�W��x'cS�J)��J�v���eNA[- �4j��E���v�ւ���`'x����W��_�n�ܠU-0��Qc[���Ug���  �/H�tz9�G
�9]m�t�}��`U�뱐�~Ӻ*�f���.<;�`�������]d�X4u�=2$���2|�K`���J�;��9`_��VdZ�i�޷��J(f�nN%;H�&e���NaS����|�")�ՠƟ4��T�;X9<�u�O��R�u��/������Uϓ?_��:�p�Xp��[�W�^�acػ�X�]V��~1�o�5�y�����w�}�f��b�^����Ph�y��Ь��>;�^^f��ҫ緐�?
C���{];"Iɐ�xiQ3�8@�s���ûo��j�.x�m惥��y�}��:[=�CL��Or���8�,gz�%5����bp�!h�<������X�
kS%��V��<K�Y��c�u���;������O��]x����Cjw�+�K	�D���/�QA<��}X�Q`"���c^C��Ә���5U��3+g�G,���f<U��+rn뗔݃�МU򪕡s��^�v#,#J��׏#"�4��[#`L���+u}�f��$a�<�a��w��,a� �@ET4s�e���*@hj�
@h�M�O�l��zZC�)l�;�TӶ�^�,hz� ���㫡�j�=�^:��^*<{
������1�u] ��%�f�������op�X�7M����a�ir`����^�ʇgqm�w/n*��Y�!�N�6�d����d��@�2�!C�0R(�q��t�K@I��Ϛ��h!�n�r;1��b��	*�1E�������T��o[���A��ޠ��u���2��ܑ�����Z~�hH:^9º
3�u�,E��h^vO9R�Jn��c��?��o���H![����֛RGO�[��oJg�����oBG��>�ߨ��0�3x����k�xj�N{���r�@�-�aT�b[��r`�'���ٸ/�s H��oN:��kE *=�~dՑy
��x]Tp��gx��Gr-яo<��_,q�T�����,�V��7�%7^�ƶM�KknVAd�f��1(��l��~b�6L��C+&��c�	�j.b��7�!��|��)3J�@�T��d�LAJ<=�����Dd�T�w^^����󦼒K���g/<w4jS�$t����9ǘ���$�݀vZ]&ds�(�4���?\˅5��=t|�Y�3�5����u�qA�P�Q�6�~QH�30=������1���m��_r�ǟ6 *x����~�>ߓ�]0u��ZVa����IUN�+�U3�
�'?:F|||���sX�ΐ#٦�v	����p#$U89��r��a̙騅����2䲫`u�F�_�Aߒ����<�X����[Y�}P9�_iL�$3kDk�RH�A����>p/}�!
ȸ�&�΍�E������w�@>G��GVZ�Y{��V��ޥ���_�i��,�Q}ݧ+���44@Y=�۰�z�V��>�����k��##Ҧ*���}�v%Q��K�5�ZxM���������x ��wB��p�v��"z���
^dH�
��`j�t�v7T��'��甪��t;;m3�H�Q@�Ă�4Rm)�~�<&��?R���ӽU�� ��������a�P��o��4��Ӕ`Q;����c���8`�G	���@M7!����3 L	2̓V}�h�۬��V%��<���7ch)�e����8S�βֆ��
�Z��	1x����WW�� ��
Zz��\4Ҍu%t���.甼�K��Ѥ�/n0���(�^�N�2D~��M3�q��,y�)�c:n���F�6���eN� ��p�8-�I�-i=qWX�	
Z����z[�A�����r3��O��
`�c�a�\�~�h�C�2�/'�.�NX���9'V'+�K����.�v�X>!3�2j�dp8��`����B��P��,J���f
[Y�L#�ᢰ�`Xv"�:�c5 ��e����>��w�0Z��|ei�E�`O��qT���u��"_]�=ZM�.�ذ�2��\�`�^�ྎ�Gf���7��l�o�M4�� ȴi
�z	��t����|����ަ~�vWWCNtC�N[���{�U��	��[�
^��\���a���G��K�㟸�a�D��W��~���xo��@P�#�RQ�|R�#�n,g���0���\���ԬNl��,A�z�k�޽,-��,�/.��h|y�M*�
հ�a-�-�쓻`�^�,���;�8/WP���(As2�Aq+�[A���^��&�|� :��x�Ī�Gº��{e.�`�0�݂��z�A��<[��M�Z�`M�G�.XzGڊ>
�c�����K%�$Ô��vf/�����?�y������Ѿ���X9R1~Wx�j�p�M>�13����|��՗��Pv�K˪ǰ����j�ӈ�u�;'l�K+Ҷ����d)�$=Q��k�y �~S�a�_��"'*�m(|8�/�V+�l�������4C��h�7�Э�y������odےZfkA\����wH/t)����6��I=��vp� ���:P|;�0�.,�݉f�uXﺸ_�J���q�MgQ��i���:Пv����L�I�f�^�r��G�|f[X�w��n���H������D2��o�q���8j%�֤%63%=6�v�;���2����|�כ&��x�&�||n#&�K_(	��|�y�+��?��5"΢=F��?:�ef}�4s�ygvH�3p���|���h�Z�����s�?��N�z���QЪ��K0j�/����r��G�<f��]'iAւ_}�|×>GA�u�1h������/�U���V���H}�)���7����:��tƇ�$��n6��
����.C��cXtޅ
�f�H���h˚j�7Ո6纏��j2ɯ��j�T������3�V�ċ�U��#MP������֣�S��U��[��k[��P�8��V�Z�G��7t�E�ʗ>J�~�pd*x�CDT=�Ѳh>�����Bz[�D>7�ʇ���
y-���Ϩ�C�;�5����`G �c�`���A��������
W�B��6���=�Ǻj��S{瑭��폳��������D��#l'^$���*ϙ�1iAM�
:��3ɹ�S.�l!��V�W�� 'i��dD�w�*p}�c���Aj}�q�?���V!�!O�i�S���f��	���I�&{>0�g��U{������[v�aZ?��ƈg6��W$fN�H.����]�:�23M*hެz�#��ْ�V�G�����ں,4U��!W��s\��ô@sߟW7�����GV�=��m�t(OC~�D�i����"���c�G�VfI�$7*�g �UG����e �_���Hi�ɠX�P��=[7P�Z�&������:�� ��!�&~���'�F�j~�f���r-�3���g���<�Z!!��}v�ģ|����L�j�y$�T1V�i;P|��u�*<��-��-���<K6�J�֛u�hu�|`���
'��lפ� ��.�����K-��+;��IE�hN!��\��<�=m<������x�Bc�j��V��}HDi�ؑހ��7��3r+r�T�#�5Iw�Om�XY��!9�ܒ��L
��=� NQ�K��Ȫ�V��ֆ��.XM���Tz��.v��"�׿VL�e/���}<���qH���kH��`�g�]�d�����Ԧv�c/ë�֌�q*��{1o�`帖j���E�-s8�k���"��Ú�{�a��>������k}I3��aLe��k����������G��S���?��̤Tn�+n��l!��=t��(*M��'G��ۜ���|7%�"p�Rrm=������]����y�k�z��6/6�h�q�$|˒�]��v;.hk�os*�a�K(�	��oM��� �	}
^�w'U��̀�dA+�$f8?w?��%O\h/k��#�����Ҋ!�#[M�pX�6����&O�%̴�X�8���Y��ϵ��rM&PW���c�~�ȇ�:�A�`<L�=���P39F�qU𘛆�=�c[�0l�Cv�ap�_�$��H�����5�L��  H���"v��Y�V)b�xi%湺��x��d0t��Y0g��2��kcյQ@����Cߘ=�fa[�X���(�h>���%n��>*���:����Z9G��z�=;(vB��@��W�Bi��ʥ�R%
�;@VNU\�3��߭u|יdI.��6�6�h8솽���(�R�#��5Q�l5�y�w`�,�#��������s���X��c9x�Z����=�Ѻ�RG��m����SJB��aj�4��k�v��U�u�D���(���&����j��P��R��?X�	ܪ�@����N�w:��ܧV�������$�9�6#�Ɔc6@M��:5�q/�1A`Kq��>w`������!� UV��c�)��a���k@�C��&��U���!X�X'A��#h+dM�����|�����m� ��^+�V�yI~��
��ɲm�#�����S�M�*��Ӭ{�a'h�����{_!7[��3#�l�I�ؙ�A9Cq��[q٪�)}�8h�^�EIDHVV�;������췪NnXT��o��D�R��]�U��bG�#�z�&�C��|Pb�8�[��M�8@�ix���ۍ�݋��&Jpu��J��T�蘵S-����d�7es��N,��jK"?5��|\�!�
3�z���~��gL�P�EcP�>\!b��MYD��ph`n:���tN�w�,;4�����o9�k�S^�}\���E��l�[v�gE�oϚA�ʪ9��g~0[ëbF��]ѻ.���S+0}�Pn&�JF��� ���!�!�C+%�A=��k� `l�}�I�4{�T Z��}d��k-J����5{:,�#}�$E'y����Ǟ��/8��C$퍬����;n�>h٢(i�
�i|n K㐡�s@Tvjn��V;�qplG��áC��cIu��	�g��2��|����\>�$PG�-N4gQ���XD��<Ą���ʎ�Ab��%t��Y���h��YЀ����%v�ʹA���7����\��f�<���� `� VS	}Ֆ����~l<�b��ADD3v�j�j�V�� ��p�f��n{~됡Ҥ�̱��79\\���#�1���$E�xiS�v1��pͯ<�,�X�Wt�����HFQDM6�K*K�c�4�c��l� m�Ϛ������I+t�o��ʶ����܉��L/^�ݲ�=Q\��"H}&��E�+�Ӛ&H �M�;�]��UmĠ��9�����>�:��
�՟��$��|]J�o1RG"S���u���^��|��V�Vv鞙o��	NC]�0y�w|�^H	'-�q��C R�wE�՚���E䔠;k�&t�4xxw�������� ����Yv'~.O�#4��Z��<&J���j`�˖h<H&����R\�%�g�n/t̚��ȍ+��gy%I���@�H�|P��^�+FX�`<Ϧ���Pn���Hv�4 �W���h#̢�+˽4#aih�*R���ZU%j�&��w)A~�S��<�pw����A�#��+g˓$��3䠡@�g�{�&���'�j<6ж�2}Ը�����b�y/}�mh�ݡ�0��`�<6���Jjj��?L����)�!�%z?��^Q�������W�U�M�ʹt�3pޛ�S��̌�������0�,����_6�d~
��ϛ�d"G�C��x�����`���*��D��)d�����^n���c�0Q�Ȧk�;\�0�]g������u��̖����c�S�������`'�m�(�yi��լ���ÍY1�4�� �o�	��`�2#�Q�:��M���<�~A�)��/ESb��X�5s ��Kj�I'���s(��#��"k�%C{��PR�B��^ڌ-[����s��� Q���GG��+v�Vɇ'Gn�à�γ��ؐEf�����4��7��}k~3#�ަ�ޝ��}G������aG���OCV�)h{�;d�9Y��ڎD���y��5;�~�k�!�����t��`�KN��k��9fKT@%�ύ|����������86u�I��Gv�!Z�!9XjˮH=?����@E�����j�ƾ����|�=�`^�4eA
��BO��')ߋ�f`�pX��^�3�jy����5����$@��uy�K��j9iA(WqN��|���t|��CG.�Xvk�Ճ�b�Ƒ�w��x4�gl��Yt1-	��ٗ Y�i�*��%OU���߽�߫ۜ����E����p�L�c�%>�kdB��W<c��4�cu�Ҝ!:��e&⤫�CxVI�8E���T]+c��pXOJ�c�w.�)0j��6��4��
�'Dk+p�M����6���dp���F:=�
:qY�=Z��ԪuP�Z{�H��f-%�����fs���w҇��x��2O	����l�oq�i�^�G����C�!<wA�;�yX�Jn����)����p �����S �����=JH����P��jq_t�]+��\�nTv��,�@������O˭�9ORk�4$�,���4C�(���3���[���0�վ���H�r]2y�Z*����;�a5���T������ݞ�_����%z��`M�G7 �Wf�P����er��[�p�[@����_f�,7J�`vV:�����m��9#�W���/���YZ�+��������m2$2]V��W�'�vʗn'�ykKq��@�w\݁J��Ϗ�m�5���
d[A�w��piz5ʼ<���e	Ād�Q9�k�������γ�;ѳБ�᫢�Se���N�F��^�D6{�
�rǖ�L���OV��
nq��e��0Γm�G
Ι:�3�H�>�knrGO���WC�6	JƆm�\�F.	>ܑ�XJڙ��Wp�H[��_�>;3(��ݰ�CB��<�A�l@�76
�wǪ]]����A\Iok�Ƈ$ᆝ��?Y�t(�uS\�����\�	�Sn�'hb�M<������^K�uA�9�˚�R�ӿ��~*Qh������K
_Cy�B���Q����m2�.I��?���g��I���3~��y!����_�;��x*/�SՖ�z�n[}�y�#1"EC�i�Es#e��uh�F���-���.Jz;���p[��2|bk�(�^w�.J����v׊N���p�%�H���JՍ2�<�B�u��&�I}��5Re����hPb�X�N���Ty�Թ��#�[R9p�k-ēUFu�Ҽu1�T��i^l;X�����E�:�^T�.�P��։Iѡ\ޜkd�/�G�Ə���%�ts����?���Ks��m�\�xz����&����!aQ�^k8p�@ʨ�Nc2}�Nf�����u��|;�6Y��z�2��;d�v;[�"���Yі	��VK[���7)L�����D��ų�a��x;e6\�?�١����@��H � ��3e�͆I-���]��O�H&�MZ����V������/\�����ɍ'����o��́�~�����1S+���1�7g�K5�d������.!]�ߚ��}�k��Y��J:j�W����&���=x��\b�s[K��F#�6����;m�6ڳ�$)��й�X�#��Wp��f���t�\��	�yh�Q��e}�yv>uZ-Cw)����-\�n�q(�od[-/ufo �M��)������'���2���gsr�wN
_�^pKF^;�y���V[Y���~�y#=�/��k��Xg8�&a�Ŝ�?�K8����ĭ�և����<,��<���;u��1N�N�����s�E\�Z��>��Pi]3T	M�91�"h����Hd;�c4���>>C6���7�K0z~B1�U�R%-w����r��[�PUmE�Q�lC�MRg?�mt����{��\-�1vh1��[�Ha�?Ś�Ί�GG�.C�W�:jpH�#/_h��E���b}��_KM�ߤK�P�x�h��CB��\c�� �g�UrU)����e�8�ly�գ���Y�AU�����Uq�%+.��*몔t�+���rFx+ �1='1#"�6�!�/�#\>I�?ozģ�U�|Rv�YC��߬G�WXR�_���u�Hz�Z�
�X�h�{P5�U�ĦڈK��\�6f?�p��vp��u���{��8%��*-���~gi�J�m30f+@u��!���
W���u��ا�;�%�z�ǻuI�;
Ъ���xiJO�u�9b��]�a�òev!~�֥�ó[��*�Qy��j*�oe�밉��Yz,	�^�ͼ���߮l�`��<�5n��u0��q��r�XZٞp����~fmIF�/��^�n�y�*Y���El�)��,#O���ޜU�>��r_�{b?g�-�Q>́��6I����k�bu�F���*��ׅ�?�xW 6��ګ1��
N∢R��I��+���)Z��>?".Ñ*������G<C��{Ҹ*������%;K��IP��L>S̨�	�d� �a�/F��"�[�ӕٍT�2ˢ@�o?��%�u��c�^�񗞲�zOlĔ��[�|ccGh=�㧝bP2	�6�F\��)��>ҿ�M'Ҕ�2%��)��=����}�3�G&!�9f�]�a88;���-��B�������pp�:^�5Y0����v���aS�P�w�!��([p�Ύ��H[����w��8q8.5��?���S��X.�:�n��y��}��H�u4"�ɴŰ�bP�̠�J�^�[��)E�׉��`
���4�e�,�~;�M*��*�D��qO���5�!R����a��qeb�R�+���.%wq�g;!oiC�ۤ�6{GǠw �(�Y���f�~�������E=�p���c�m��ۈ���ד���9"�5c��Ha$���rpi��7\�x��t�ߞ�ۑ�V�s��6�6�b��k���;��N"�����L�$z�2E6KHwO���Zґ�j��N5��U:nq��z������la����U�K��!�rq��7�p���tS���Ti2��J7~�85U��H]N�'|Te����T��γ�r`Q(Os$G�����qi�LK{}��|����a�L-"�l�������������xڳ�fY9 :��Yv�f)�QB�F����+_�g�\�RP�
Иmh����CB2y���|�!Y�)��KQ̎7���Z���ZmzFN����k��}p��"�M����1�� ��T�C���/�!� K�ێ&�
��RWĕ���
f��{zEC�C��֨��j~�{�c��Mvވ�@�\̠��咰�*/��/��FE�lq
f���������ٖ�~YN�����WD�������jr��M38��j������?�e���z�"�
���cSƿ�r�3\J_����7x��
@�R)���A�9d��o��֝t��AiV@=H8^��/�Xf�(�tG��x�&�r~��8o�Ӆ������_E���'��;�}�i���MԖOM65Y�~2� O�\�84��u��sC�(d-R��gy	K/���~9#8M6	b%iP��)�����>��(8;��^d�T�UJ>E�;�[X����I`�W܊�0���3Q)��B�v����ld%z%�*�1�A�R�#�6�[T��:�0/[⃔m�qb1dMY�Y*��k���l���g�������v؄���Y��G�o5�h�+~L�G�'(��u�-��^=��B��"�R�Fl2i+�_
tts��:�s�y��1�?��o
�fgޚ�^��D:�4�˞`���p�뵃�KoM��60Ӈ�A3`�b��>�p����J.�+��Q�2���a�;�7��c�%"#kD8Y&R=T�#}��X1�$�nw��TI9�w��uM�-I��0;�4�B��.|+�Q�?dT`���Z��x�A�P�<p�3���F��1yr�1I9�Fr)��#0�N%t���_� ��J޲�!�B {A �r|��N[�kAA�� ��R..6�Lt�C$ �[;r�;�%M\�s�-PΙ��YS�%�+�0��'��s� �Hn��%�ft}��pȾ�����H���b*sSr��'�C�Zݻ'��0��l"ˏ/�|�eqW��8A^UlLh#���	���Jq���' ��+֐��m������Wl�HJD�+۲�TZ{ܨjS��5��h)�88���V1�?��B���'~���ɍA1hpV0���S�ho`;ڈ\��'^b7A�΅���M1���^���,��J��%D1C��*�g��/q�NN:M2zQc5�r�`�<��=�'_
��SX$p"�7�#	f#��(Ys����#Fp�6��:���5��M���
�3|_��W�S�1���BSн�;��+	+-�Hz�}�*�8?y�Q玖3����R�5Cyi�D��!���ն�Z��Ԟ���{�Z#�dq�u �����Ր������<��� �o�R�>RJI����+��i�E��d��V�4�m�����o!�7�"�ر��ˎ��+T�|K���H7�V9�k�%�:!�v^�����xQ��XŌ��\m�d��*�,������}�?������V����-4��	0�U�H\�.#�S&cn�@�v{v�o��)�S��s��k���B����m�=�\QG������W�il*F3���� 6F���xh�Qe��l���ь8�HJΙ�I�s�"�ܐՅ�߳�w�fX�?�ͥ3�c9K��ݚ_�ڙ�p��A(���qA�d�=2�rC��[�%6+��'��h�2�'����Cs�ĸ7�N+D�
��h�Zm���O ��F�˕�b�5m�7�ۏ~���Z�߈���.�x�x]Z��S�Қ[Te.����(RR	i{������aɪ6�Nd�E)i�R�&�VP<n�wd�:�����4g��{��{l�ς-b�u�_�\��R���r�֤2�$�")'�Fpoρ�]�͕CU�y*�b6Iˌ(�޲�Z;#�+�[i��K��|���X�e}���%/U�@ 9._�N�cWS�b������aA lsѩ�����Ǔ���xࢎy*���.{��	���!�m׺��nP�����Fy��+3��3d���Fmr��xz��yz�x�9ϖ�q.:�q����O	 {�?"h��f�����V{�V�0��S��~Do�?�>��pf�yF_��ףM�(g]X��P� ��2��%uZ��=�Uu��n�-�=?��'�\T�1�a#��sM>��6H�z-�>�ͿG���P�tw.YbӘ����T�9:�^)eRO�{8��~�y?4H�E��WX����VV��A��Ε�'�����=C6�F��
� �d�j����]%�~��-�1�������#èE]����Z�q��q[_��v�����SKM�Pm�5�zZ�j�����Sv�F���9U?��a=B�o��g��!ݺGzWg�� (�SM{u��k~��&s�bu ��OA�ow'���욭7J鼦��m@�J��>bM;�����8%��؏�h����*�X�8�j��T�uR`�bu�G/L}`��|~�S��R&��г7y�ܡ@��(��0w�[��%��Ɵ��vf$jH�b�%'�,2�W$��44_R�CFԉ��|n�Vy�@Z��
~ъt5�֜#�d@�{ŵ,�
��4�8hqX�OTv�q�rƟc|��W�HCU�h��'���Z�Ј�AQ3-�����~��wF6Ih�QB�O���Z5.W�J�eKOUq���%�)oT�pB��*�pŕ��,�8h�/��	��=b�j#�"Qn��;)п��Z��~�\��Q�K�n�U�L�A	�R�
�:��!B�>t�ދ�.A�7��ȫ%���8.p�`
�{�4B��{�5Z��3dּpń��L-�.2x�P�S���q���f��_S�iځأ�v �A�h�@�bhm�Ju��������w�E�pE8_��^����%JP@�[i�k��~"A"A�eǞ	���H��.F�n��b+��#�� s�ˇ��ࠐ�W)&}��z�Ҍ��Ҏ�a����!3��d�؛#�oP@�$��:wc��ܦ�:����Q���!PTP�lT��"�?��݉*��m����"�n��0q�M��c�ه~ȡ?�h��⦾�8�m�p��UX+��S�?������"m��t�6��{��Y�_�=�̮ߜst��P�!^�x��L���;U���������1GȓB J�*r�ða�ӯ'�SU����P�l�C�6Q:����� E+?��b�6T�+Hͧ�f*�MڠyAjEE�E ��UAE~o����㭠�g�>hb豓��]�	S�� ������N#"�:�����3�V���et������'��d"L)�TJ�NB������j73���
㻑��	�B�/����1��~0ⱽ�-�#ѽ& �s%�r�B_@�����?��,˂��V������BۜȐ���	i����gU��ʵ��؈�h@�x�����7ȯk�ǡ�
��z��_���1��՝���u����+$hU)f���|n;2mY����[`�]L3�@�?mU�%�C|4 |,��S�k��Q�l�U�NP��E����P���z������Ϭ:,{��C��F��o�H�e�0��T�D��&���q�@��T��#��Nn��� ���%�h����OW�I����~�#�W.�Ӄ�q0�GDƜ�R�8�#Ÿ���+te<peɽ�1|�g�j�,C�/��6���G^2Wl?�����ϡ�X�W����h�kw��u	�{���%w���M3R�
9�9����;�V�L���+C6����g������/�5�SCB@���\��,�|`UƔ%(г-o+bl����L��O� S����=��6��`�jëeK|*��l�D�u�{9�0Z!V��ݲi8���T���	*� ���͉� ^fZ0B����ʅ�	Ј}��2�;��-�Bn��lu� G�V�.�E�j�"���ƕ��L|U�t�_ѥ.�̰�*:��[P��m�E��ĖĈ������V/@�7�#ı��̃X�8/��#�nhN%ץ�dl)~�05�f�g@��j�	�����!\�ʎ��.vk�"M ��JH>O�}b�y�"��������!!�eT�>����L��x�i��3a���X]_[om����uE�� ��j�2��B\Va����P$ >�`P�O�����3�g��fsCTڗ��!f7m��H�?��ߵ��G߹��R��B7���_-�?1(��Ȑ�3�`ۊ����m+��e- 0��π5�by��<	b�����ܣ�Ou-��~��|/�MY����F�B�!��Ȉ[S4l�h�h�a�y[SS5F ��[m��-67� ������x������ݣ4S��.2S��qP6<f���o؀.�(`���4h�޳ 1�ԭ/X�G��z�k̍��Z#`��F8�;e�S���%Q�Z�rK'���- ��Zܙ��,QE���Y��W���aN��{��
�`p�̻�KU�^@�@U��mc�����ݿ�gj�e1��� ]� ��:U����.\eW����s�<u�t��4N�Ha\���*�KY�*sw�4J�#�e���=��3�����?�Z��(���ݧ���$)���9D�%���yt�N����W��=Q�dd.n[�t�p�V-�Xu��>�S������-n�!���x,�m�Q����Q�"tC���) ������)��h��[\:�wu��1\8:J��}���=�y3����I�0Zu0[��8|�G�$Ֆ��5W�B��bj%ܺtXMH��S����m/�*����YhMk�KO�����pe�[S4��zB]&�O3i�,��Ok�����4aM�x�#��`�����
<76;����p��K�U&f��\M�"U�|��з����;ɸ���+����X3�ʣ���1K7q4�~pE�є!���U�A�-Γ1iD��cm���h>J��=	.�l�b��*~��˃&ߩZ>UmÎ���%Or9%������*�����_�D��CK�A-����U����!��f��aL����˽O�UA�z8�&�P���ϯpd�Î}N��(`C1b���p10\�;�u�9���?#7�����2���a�RD�\�(�ވ3��y�c&>�Sz�p��O�V����n�8�ޤN�"�
��B�Xe�'Ǚ�3� j�j%kw�/�v��G�\�(�aI�����u�XE]n.j��Q<OW�\�˥�b�������P���a�����أ����mQ��ә��ع��#;��l�LN�]�)��ZΡ��ǿw61�|,U����1$컦B��ッ�s}V����&ͤY�FN<@���o�Rp�Y3h���	/ٚF��@<)�т���D�0��&+��χ����aW"V���+Ή?w����c{'K��L�����B���H	[�t�$�t�D	pm�8�%��]�߮��+W��mo���M��8�SZt�3���̠Fd
���?��Ҷ��S�ԣ��<��"BHHН=12J��.��V3�Y�n���?`�$�s�{n�y׻%�Oc�)>�*�<�\���~�!�p���w�z-���Y�~��=mf�p��ċ�ʏ;\���_:��"&�5l�i�9�A��(-X�e�He�$α������2h,�U�nʸ���(󨇥�>��5�0g�ܿ&���C:/nW,��W��5�ehЯ�C���3���t�����x҉���0�f�a]g�ց� �0��G������X�����Iyx}���Y{s̔�����犻�pX7r�'�aU^�Ē�������UM9�((���e�II��U�>�o�/���
h~�<��񳦮���7̷�$I����eУ�Z�-�'P�$`��0=���a-��q����3�G �Β�]~Wyi���x���4��X����1��JSH�4�(�f{$f���'���E�Hm. �����p@�i��?*�#�Uq��\8e�xo�����ar�$�K�G��p�h���]I{1v��T��XA�'h׊�ēE���6:��8�H�j�����"��4[]�	��Ұ����Ui]�q3`a��j����@��̞����[��N2 �'���˞���\('�O�"�����~=��>f7���>�`���pS1&c���ՕÕL�-d���Z�^���E�3��w:I;ے�]0�@�7�+�N�
�;r�@c`n�޷�Ѭ�;[�n���v4���_qÈ2��7�]$��e��t+OIZC�A�@�oE���N~��
�pқ�	gpK#.�&[��C�*Vop8�x�P�@��e
���g6�oe�3	�G�����s�hV�t��/aO����p�E��+s~��ľ���\�~�����S'�mVlk��� L����̹��wml)�ZF�I�����!ʶ�#��?�2Z����/
�w�||j;ȉ����'��].!�_]���-~��$�ϴ�I�Ǹ8�?��ߐݐ!G����̴M6}����RQ+ �|�d��/�K�-l���Yo��'�z�w�3:�a�ޜ���2�˖�������P��Ԕ��l�;��T��	�.���F��,i��xY�Ld��S� �}����J�-5��;����Ko�%��U}_#�����'�fm!�ds�K�P�}�b)A��g4�^�)Hvs9�MZ+�0�����p�*�����B����~�X�[�;e��ʡ��G��#`�8�5��AyIz�x�YIj11��`�֋���eYt��RWU9��I��/�@�pX�$������J�|P]=��?�6߽A���P"���G��ey�	,W�= R8F~���� ��y������Ǟ2"f��m�X�#F�ڽ��Q�ꣴ��[(�vݩ3�1��nc�Kzv�$1e�( �a�X�w�2�^��\��$s_�g^胢֐�~"ހ�S����aW�
y+� |]���%{T���h_x��x'��{�¡���a�/���{N�����c-�{	S��yW|`����$�)����5��`��<�f��}y�/NEU�]!G��3�~qF�D�h��O&�#��i�	���Ͷ"%C� .��4��{Z�pC��o�����k��� ;8
!(�;s}�&s�����a���S	r/]�Q�j��4M]]|��XT�?\�o]ue����؀>���JY���� ��"���PЮvi*�a�=�_�L��>�#bI��Q'
�,�|�yB������PQ��s��#�+E����*fM�d媚��tS�<��HH.������Ćy��$~ڸ	J*����Pƿ�2�̽�q7N���\~E^ޭVe����% �\bt�@R�]�,qϻ��i����a������a2�5� Rd�(Z���Zx�b�p�>��m���7I���C�����\��p[�$�@�����&g`���x֤��0�ܭ�	Q��̮��cS7hQ[������K_(ퟱ�$ƈ{|n?�$�M�;���	& �d��\c��_�>����\?�;#~�f��	�e 0YwT�^�ۗLCxn!A��#�3s����O֝�#F��2�M�>���ajʽ'���,; �e��-�}z\�,'.�ZPlh�~P��bx�. �oS��m�R����A���L'CrD�t"���{E�����R�s<�Mxp�����Ed�!���������D��蝵���$�5e?�g\}������"�/�H�,P�:9�{n�w�_Xu{��#q�,����<�����u�P����ఆ?s�p�/	��Xº�Q��ѩ�IG��編�\`��}fh�E��/A�"DV'�Y!ｭ�
yt�@<+���D[�qcd�'�"�I�n	9��oV��W�ЗJ�}��@��2s����l�G�i.�笓xW@�`�vc�}�biU|�K�/N ��j�����>Z:�����?�PI��:B�*�<��M�؇�'��,~>/�����
������&��<�٬Q�ܭ7�%h
�u·od�� +:�̋
a���,j �'B�{�ϑ��BQ,����v)�� � �^ �~��lİ���Vf��-J~A����L]u@T��vX0 �DRR�t¡$�K�Nghp�I���J�J9JI+ �R�1���	�?��}���|���n����Rʺ�B���a]`d�9W�l�9����-�qr��DQG���_~�oXx��(c��%ٗ,BӢ�vP�� �/�f�a�#��h=���#>7�|�>�l�/D���{KvP����L
�RI��[d���bo���U�D~e.��Zwy؞�{�A�����;H�H:N�؝� ��-Y��62Ia��Qu���ٜ�t'�)�	���S?Q/b<���T��WV`����_�L�U�m�r�4�˕ %��<<3֩�K�w+g�s�Q�?A~
�~j��؂��&!X��.n̘��ӿ�X�9q�m�� 	������Q�W6�l�H����w��jNk�QO�h�PXe(B���/V��B����P&���Ax���{�*(������s���������!g`�S��q��s���%1¯'�	a_,8�Hm����"4�Y߷-m;/�����R�������C��y.�D���Y�?�E����P�؂����|*2g~j�2b����)�P�m[�t�0DFE�';a�����U00���o�9�a�M\�YS�&�-�C���Dq^~�/�vp��!%䍬����C(#ť��3C5@c�;������KDo�,9��%�_����Im�E �/�1%��-W���|�a����vh��~y\�U,���|�k�E��ge�R�D�Ll�;�5�j��֭�>��0��-�����:}?!]�X����e���6� �Oӌ���+�?3���C�ߞ��S��3�J`�z��D���z�?�L�L/��-�$��^͌[�/��c0�Y�U	f�	�/��o��bo;/o(���D��+�Fj�OR��0����c��*?��f����� �Q9b�\�C1��l��wz�f4���!0�QN�j*�:�s���"̤��S헛SR:��9��}Z�&��bA�i�$��m�W�4��q�VޡKꖗ@�]�F����������Ì�N	X�w��cCܠ���τk:��8�5TTOgf21n*]
��7��6��V9�BUM_�t��kG���>��RX9�8�Q�Usv���[�Ч8s��i0���A�:�~��߲��B<�[�g�Ys�O!W�Z�� !�/�
)P��A\C.mO���fec�3�ÿ$��2����Rj1�&�u<� ���R�&��	3�iĖ*��p�� M.��)K{����ɴ�M��p�?L������+On�����ު
���t�;�A>wД����"�@�/'W��*�����h$�{؟V���$�gc�~������"�Tf��b6�|�,��@�'y�����V�+8�u`�C`߃0O8Y2,�U��"`����ŗ�>_֍�Dt?
$��v�"�/��oA��&
f_�8��H<�ޝ�fq��j���U`��F_�Z�i־T5����wP�S���/�O��ւ��a�~�1�R�����˺^��=�կs9$#r��_�@t�W3n�J��̏�����g__8��t��{~&&��"ࣗ��O��6�)W?�P��\���G���G�ɑ;��
��?n�ɱ��p֛(J~so�S��vn�9�
8��!'��!=�Hz�*B�n�jt�*pΏ�'Y�9a*)A�o��u	oPoh�a���"��KT�;�x�=v� ���X����9�cf͌,5$�������K���/~�O�SL�|��]�	��	O�[_�xs��\37�(hH��܁�vv�@�����p���W���7 ��9"����FO�Tn^�[�m���~���N���'�,.Uq�1v���u���;M�Ф7�l8�ʨi���A���7`!q6G2�%�4G�6qW�m����~���R@$�=ZZ�Դ_�Z�<�.鸀� 
L�y8vX1����<q���Nz#羏��da&)�~�&��O���{.}l	�WaFP	��p������iPM��C%�O`�p���n_�[Ҍ�$x|��Y�uj��bm���ė:&��g� ty=$<��S�LlnB^��&2��Oc3��������t�_�]H�D`0QY���gc��ܺ���́� �X����$8l;C���@3����
Ǻ���Ӽ�4~�ơ1*%W��YR� S�������3e�����4B���o-�O5���
R�.9^	���5N	��M�~���WYW��|��c0V̚vi���$v���#�M|��Lv���7�X'ر�ڂ��s- @��]��~F��N4���W���0�IY|`���O�m� ɾ��\`�M�`l ���`G
�[u��+�B3�q͌ǥ�g�r{���EL9�&���K�F�rr?+mKmC�(�OgKjAH�\�5�>�D���$NJ��]3
�6i�6�mA4.ǟOs�q�&*��ۀ<^q�>�yJ �;ks�b7Wx�p�� ��/�М0@��@���$%t����uzv��7<�R_(�+��H�Rf{2(x#�b]�rNKJq��W�D��a~����]+��!�Rc��\��}��`��X��b�Y50ޠl�D\��b�#��%6�|~�W�W�P�^
:�� (K���������_4��ȬK]�řH�1�1ߛ�<3:~:S���!^p�e���1�6��r�b�?��$�ucB�d#	��Ƴ��1�3��fu>���D"���wnճA>�d�d7(r��y��e���ݏ��Zy�oH����*�Siߐ_f�T�����?{Fw��D�,;�]Rm,E ����b�O�ϕ�,m	nঌ� �sx86�{� ���#.�-=ҩ�о�I�+��aﺤ�k{�����@�c���fu�a�?��P�en����jOpM��=���A&���m�I	@�a2������Wx�_�������`����g��	�U�_�IQ����,��P�'���r] ~��#!�։��[E��dn�?��IP�����_�����J15�ҳ}�OP�1��_�fr!J� a�Oi��ro�R�8|���y�O�&�������j���l�!����3��G��U���w�M#@�	���m�L�O=���)Yۜe�Hztu"-��>Ōq�m�)t�K�t 9�֖~�Õ�4���.7Y��)�Z�2�><�wm�v� �i蚍�7_m_XW��U|\Nx���9A��2�}�f��)$��?���X!���G|��������ng٠%�<�[���W�V�ߑ��^��)6�}�L[��
yYy���`6����"�[��
ӛ���O��5R��P� =�Dr�|��'6e��,߰�?�<�ݲ�~C�=+�N���_
��Z1#̓���_���(��.�Cϱ�^S:����G�Խ}8�q�-���!2(hq�̄�y���qi�@�S�Di���`����߿�x�K�p�8��}����OϿ�L�ކpp�i��2
ZR�]=zUwh�nnM��;Es/һ�4�
ή��p!>�䗻��"���w���R�,�A����~��i��No����S^�Z+f��I�C
�qT֘^^9���*�t	`[; '��s�g�hx��,u8t�9�0u���_���=p�}Ph��`����d�Z�jY]H\XuR�da�����#�u���ƥХ���������BЍO�����E�K�ߗY{���`���[G����eZe��S��%���y�-���&�,���ss�=��gC�!�ҭ�j��8�H��g����F�9�R��و�i	�<��g��h��oIIP~h]�B")�����b���1���I�b����s�}�2��b<��IV�;MBc��.��)s��с�\=S���b����́m;�)���'����u�������Z�c�I6�!1b�Z鶲��H$�J�ѯ�cV�eĶ��S�r`da#���-�v��$0��Xr�W�N��NIf.�:�̼�Xd����!{^��V.y{��6O|T �;��l^�,e��]g��1������n���y�����|��C���	�W��W�9�����U�b�����p��
����d���Њ��Ί"b��G�pq������n�3%�D��zMI�
cZ�H\�$��Չ��b��EͨS�	��5BYZ�Z�*u��U���2��ᴕ	���O{�i�S�h)�p0sCG�����𩍚q�9l�%C9�&n|sd�_��$�:+ځ�eo�D|I\JQe�&7|�Z��t�0	���0y��і�.� �=�}���LY�/xx�����{�A��Uj�\:5�w�V:(�x�LW���|�7�-d���{�/�Pu���$��6�b��b.d�C�ӣnb�U����}%�*�5���[�0Ã{��b��,޲�v~:`��a]��W�J�Kѵ-�0/ר>c=�a�(e��%���qӵ7�|���O�F/F���_A��L����P�ְ����XSM��13.�,��kJ�X�=�^�Ǵ�u��`]+�N�U��\5��{Ey�,n�=w<?�E2���JK��},{��;XW���xW�����x�����Ɔ��"���v8�,�^�(�ޅ�Α)٫V��tt�V���y]>�Ar$T�$l���V=�i�����1�|C,٩3^�������V彩X�0탦����?/E�GWs����v����+ޮ�t}P������a'n� �g�z��WPH�)G���ٯ\�c������ԧ��M�#�m�B�{{�Ge"����V&��\v��6n�H2�[TZk\;��Fd��G��祐���_y���,�Y0�M{{�k&���/N�,���Okq�۩u�q�����G_
V��$1fKu�J�4�˝9����QE-o���d�, ����
��OW�/7aQn7e��O=�ն}{'(HmQ"-�`����9�Y�H⛀m٥d��Ecg�l{����Cn���˸�a��'�.րxt���� ����3BB���h�w�VHa~��YD67�F�~:���}�Q���ۂ�#"�Lqsz����������Ci�����տY�;y����-��H[I��J��N�	��&����5�c;�S�ʝ&�C�d~N��҉M��C]���z����F��0yb�i����H���s��fZ�'��1ہ�����˔��[e'h8k������z2N�(?��!��`���<�Q�MS{���[���e]��o!3��I�����c7�!��G;.�� �*�������o�MzN���2筱ԇJ�2|-�<4v+���󟌚Ǔ�ͣ�<;���'+O/ϔ0�!_H�~̶�j��n�"��6�<,��J�L Ǯ�p��V�z�D*,`FeZu� *��F~���X�I1}9y���Q�D.�V�v3���zdb�i�����f��Aj���bw�H%������.A�1��ei�.�N�Z��/�6�4aI�`/�fwV6X졬	f�ae�"�6fJ�dE�dV%�o�;v��o����e�6��n�0�̠s�IVo#��N�z����V�mm�33ҥ���^�ܕYv�ϝ;�4hB|,��o�`�#��♙i+��*[��1���s���xo�9�%�{��5
sα�h�;�Egp�[?`� |�1��|}�HJ���?���w�J5<D��:���,�����2|2�� ҾQ�$}���H}oޖO���AP��%V�Ud[)���ze�S��?k��p��=t@էp���p�>b����	��9[�؇��o\��H�(L��}�d݊��o�#�!�sc�s�����i���r��~��%�%�4eK5�z��y�EV�k<%��P�]�k�>ǧ��3�% ��� ����Ǚc��Ŷ
�	��z��M����3�� ���D���n���\)p?0\���b"���:j�_�����v7j����?5����#6k����N�z��������Ԑ�<��8
}�q{�sdax�5�^���U����jքӊaoV��Ɓ��|�<:F}=*E��=$��2�Ԓ2U��&�߱��)�$�]�I��o�A�<u�x"}�}�Q\��BtEjz�`Q�����=�օ�<���VX���w@U&�V�љ<�
��-K�ו]��؛��c�׈�;I��~0��'�z�7����B\�eҾ����Atc����S���祈��f(����u�=�1��������j.�5�}*��p��@��7��2/�o�܇t��IVla,���>��9	�w�7���|�T[mqAEk��`�T9� �%�4�X�S��\�1=�����1�@�Ȣw�T$��b;�����ň��Q>�����z5����}�����jJua"1�)9a��<��CS)S|��6��N�՚�AK��MG�d��er���|�}�e9z�ক��7��߹/$5HND*�j�I�l�Y�
��o�/S�b�^-���⸎:oU�h8�K!�|�1j���>��)��U
;��|�nm$����̣�+��*`��3����u�*m��D>�z�;�bcm������#'��u��aoR�L�M�w�/���t�}�Ƶ�݇��2�m��y�ɝ=��H�mjߍ�t)(��{|�v.�$�s��h�R����D��,�l�X��yO
�T��~�A�U��X<M���v�/W���5@�+u�
*H�@�F��U��:���P�}�t�0e�u�������o�Bg���7nSK��!� N�*O�m���I�f� 3-����5F�a�J��)�=�����񙙷�70��F�}�k�����у�E�����X�_�OO����-Ҷ��${�<0�����s� M{{�����|�T-������"?���)=��/h�kKm�S���q���n�O�طy�,9�u���d^�Ǔǃ<�\��d��9c[I�j�J�El�i������#P0�@���DRC$@�@�v�o�U��Bt��M��Ӕ��)�*՗�MK`(�6~��$Hċ9FU���A�j�Ȗ����� ��C��6y�6]��qn�N8�Z�u�fv&jɿM��V���ci*��ذ{��ٰ���M�t�I�����KΫx.��`�F����Wcp6@6%����@8�DӢ�@���?t����xO{쀿:���-���?�ȜE�������$���������J+b�F�p�8V�34UWw�c���sD��̰���� ��~/�t�+O����M�\�v�^P��]�R(���G��a�64�(n��"��t�A���$&���̹J凗���n��sq~�p�L6��8l��K�����Rڹ��2tԽ{"���V�5�y�PG] p��%P��*�]��_�tyvb%e�l2,�4�nz�J�H�����O�Ɂ�y���BS�lt{���{�W
�#�()�=B��!����k��7�	� ��϶���a^�ߓ��:��!���`[�k�o���'�㊵LÞh�j���
_u�f�	�fF����"��!dB_��X�m��M��>�i�ݲ&l�1�^�I�X}�2�2%��U:r�����'w�om}n�z��D��;�e�M��U@@s _d����͏+)�wJv������3�i� S����,�͖)��5�{��\b��*(��Sv�@��&���%�ߕ."@�.9�4.� ����I��TS�7f�v��&��xp�7��w�!�5L���Y6�O� ^��/tH]��ur�q��0ff�"�f��n��h��.x��W/�����I�>]H�TM�Z�IZ������O��nMD�8��n��K#���(w��� ��t�z�|� ���ľ��U��/m�;P�=��_���|���2�w��b���+�i�v_L���'<V��9������]�!��x��n��T�5��l�G�z��c�_���y�w�������|�}�,��!���F�L?}l��;��=c���Q��LS��W���^2�6'�M\�F(�t3A���\Վƀ?|�S���p͈D�����lI$��_������ܞ�ʌ�ݮ�#�b2�ko��{��I�қ��E��Cc�'s��n�m��`��C���I{��[r$؆g���΍Nik*f�Pg�2�g\�Ūu�x��2Ew��֎�������wԟ��V����5���nh�U���ů����ly9i�����[[&is_�g�*Wn�)��ˑ��Y��8o�g��:��Ԫ������7	=��-������f��8�����i�g���#�ә��E��F'��^~��d� 3���D�(�WTaBf-���;t�+;�x�V?Ih�����AsL�s��ڥ�/��YF^ޛ�&E�2��`��#�ڣ�o�2� �0nԔ]�U�9���k9F5�^ǚ��6[V�
�fU#�-ON_#��thY��P�EB�S�J�����dN�J�ч���=����"���Z����R���2���a�<����'��$:����bA1F+Wu��n��h;_M?�>�u%�����/ q�U��Yr�%�r��OZwȐ�#2_��C�4�3�F�[ /��E���{�wW�����F�Kx'y*�^�;sn� ]v즶\�go�	�+z�٥k���`=����_���!��N�S��{��/&�����[oR�z�.g�t��mp,���*ն��$=aA�i�wz�p�ra}G�p+=�r�V�;��V�8s��%�Ǜ��d� aS}W��m]���d�1g�;-�s��n����rH������n�PHt���`���['�nW<p����8R3A�������������4]��[i<g���T�����w�3����[11�d�}��mϒ����=5cg�2�g��*/7��$v)���"�B8\�b�+�txl�H�\�j��^�j*�]�h��eC.�� �2�Or!���f_�\�"�h�r�?Xa�����i�]�X��\/9 ���3��,
��R�<v"���a��kJ�x�&��5�UT�
ǹ��9�cQ�dݥ2��D�K��	�h�d�;���	^��KVk��>����hIx#�a:����)�m7��{-��+m!u���c�Au�		���,Nɪ�@J�`s�y9�g[��lV:�H���qj7��#���,6i��w/�*�1oU���缑�?H����x�& uK�ɗj�+?�Qƫ���=�V`�]-´N�K`�����p�6Z������	�PD��D�Z���d#-���c��eco���hM U�𬻊G�c!"B��=�_`i����xH�X���^.i:��2����*C~D�F��MO[��3@z��I������kݬ�������Y�t�>)�
ͳ����t��U�YVȭ���ο��O�>�ok�ǟ����S}U$}���`f\��s���"���[��^�8�Œ��%���eKN��l����"8�V}��Z�14e�K6���"�i&��E�<�	�6;%X&(�/Ye�4��th�P�����µ"Y��DI�p���������=z���g=n���刴hgo�5���K���9�[�9�-s��Y��P�~��"S[��cN�kI}��	R�)gU_��,^xlw^	t�T��;��_3꛳{$��:@ċ��r�{����mz6}];�6���#���5ԈW�7���4H��D'�A�=��~��&��M�T��l�4�/�~����T**�~{Xd�!�z���MR�h�k��\���	ګK�ު��*,�/b��(��'�.�b�Uz�����l�	Z���;�=U��`[?`�]8$�u�}����Bz�9��
;����})O�C�]5���5�1u7n�+�;No���>��tb떣̿��C�V�S?��6���q�Ր�� ���}r���Mኼ'q����yЄ�.��n<�6�?~,WcI���a|t��xw�]<i�Tl�(.�	4:�@�`w�v���p��=��m�r����O|��k�1>�����ȁd±E����i��@�Z��HU�ܲw�D�swγ�0�'/�uו0���s1�ʌ�>?�[m�,���	�jeM��wT��$-�G뮪×ɏq�o�
}~���0_�]���;[Kw~��V�N����%�Ծ�O'���v�d5�����R��l7'�E7�?�z�M�wG�N�В��ho���0���5�x�e����΁]c��EHºɛ�k�	���Yp��o�I�����6��ͼr2I�#�D{e�ޖr:�j�B蜜�N�i�#{��o�:���v�q� ���y������|�`W磴�U�%�?6�.���WR���C37�����sA{\@�lmR�@´+�a�?��0oVDk��.P�\�[M=K�hY����xix��y�H�R�h��s�>x�LI�f���Q�V�;h��J,@Ih��בx2�.�9JJ�j����?��G�~��2蟲y�<%�䔅/	��am��!����S��c�U�w�n�.p�\8D4�G���k�� ?������*e&�e7���_�Hz�����b�\+V�.��=UE���(������c������X�;�L�^7�|E�X�i�6���8Qf;t2(�[�T�2%2��(��w>|:ڞ��]5xZ@�� I��X-��T�����R�Ʉr���gLg���|��BW�ܪ���cP��	m��'I^y���bP&K@�t0��:����Xh�����F��ٌX�p>9�q��c�j�j�_Kŧ�u�����Kz��f�{M���'9�b���̹b�2Z'��3�:��I)�,����cE�0�-�:	.'b�`$�ѺqiZ��	\tZ{�0�r��,��Y	�+K!ǂ��L��V�%#���(§|��eo�sV�����������3��[����5���br��c����Hi4`�ד��!Z�K�%<���E�Zc=:9���}�h�c��	�l� gv��Y�e���6��-3����'���bRg8VE:���az)�����i*���z�1�:~B�)���N�6��,�i����iOc��Ͼ��E�]�w��X �qy���R:q�� k��f�0�ܣ��Xsϔ	�n�}1�����a����K���� �.K�tզ��v�۪��3dŤiK�a��ǥ%����a�5����k� 9����0�p�[L���-	@��O���2�)��1rG��a� ҂��~��
�U�'���un9B�%I��٠^K��6���÷:�	7ϖ��:�u���o<��nV��ô6k�)V>�i%�?�m�W҈�V]��ꔘu|��B'z���s�D�en�q'D�Bn���83�_���z�,��S��=�������s��sb)�M�*�x�)�E>a;�?����NU@0}&}d��.���S|�kί��
�5=�"!rv����j�<7#��x�#�D�o����7�ky��y~����rm�����x�|:R��?��Oe~r�� �I"%�2���Nx4�ѥ6DDFz��I�\����ܜg.qK!�
��3���lМ�t
���(����p��}�qbz��W��-ۛ�C���W(^t7�a%ÒW��@uC� �jo��ѐBB��4f�ƽ�����#����v�#��w�,L�֠q�{���	8AB�&�G�kl8LT���Jp�O �x�\U?�*/bK-ʪ���cD�G�|�{2����:� ��s.^�ȏ������	��m��J��*�!�S5{\7<,���zb�;<��<�0L�� ���?u�ܼ<�G��W� ��FD�8)U[��h@����۳�_v���/� T�./�$�h �z����#�?�P.�_M��]�#M�2dq�N]��{T�5��|�?Ȥ�^V[^+a"��*B�l{���ح���{�x{ ;���=�B��T��c(-����Ӿ�~	�Im<��h�q	�
Z;�L=2�be͜X�PyS]��d��!߳o�	��B�29S��𥇩[9VZ�'ۛ�I��ԯ̬�'�#"�.�k]F�8v+>�1! =l�oW˴�;Æ�G��3Omv�]EC>P��kC�xKUǠ0��x�sNZk�*����+&>3U���E�K��6�+ˑ�����p�
a����Y/�uWk������d	wqaB���AO)1�*Ջ��}�1��Ȕ�x�66�`�� w>/�I�����y��T�"XR���^e�����gJ�p���U4}L�C���8�͝�q�]	�Ұ��ؘ(�?FX?��~hV�>8Ь�@�0��A������T]W�-0��K2�� ���pA	(�����כ�F����ן��lV@��-�\��N�:>PYI#_��[��sjo�.fj�i3�Ġ���ZHPGw?zt�d ���\S��:�:*彍��۫���i$l,J�%�a�_�)B�Qf!�o�KQ�m�~0Q ��Z��DS@������!�B6��2%���+��ª�\�T:sk`ux���l�Cm�8nW����q^�b���$@Z #9��1�Yۜ���^"�پ����1��R�&W@�j~��E�M���f��<z����ˁ��h����򍊑��sɓ����א�!�ֈ����������;d���rD�-�h�$��!�l__^3r��0��z(�ʇ��>4k[�9����E��d� <br{�������2�2�TIj�Wx���V.T�r�X]t���M��<������^odߞ�~쐃|�,=�^��A�Xn�{�+#+��S��#��q@u�#��� #��A+��� 1�O#Em�W�x���t\ĈUFL����X:FX�1��D�Jq�H�FuU2ti��%�V_H�]=z���+b.���n*ׅ���8�9��P�_��O@b&4��:�+̭4�&��c�U ��E q����N]9T�m��4�Qv��UC�j�դ�!kfY�Qx�;'18�0�)^��len4��>��&�]���s#���p(7�H]�r�1m�I��Ğ�z�3b�M9�(�Պ��A_����5"VWwـ�%s��x���ݹ�Z��-����F��"_.�#�NxpЈ�x[v�B!'�yp1Nl�>hJU��}윒R�K^�����D�s����q�c��qo��-+���T/_��m���֌Nc�B�����mBL��%c�AF� �������|��^
�U,r�����(\ m���!{ӏ������'O9X�����]�z���ݙg��{|����$�I�S��D�� �a�ནGK��'��-��3���8_yEp��3�/��q��Bg-�9KL,��>�O�T�l�+���g��l)g�$U�}��rL@�F~L%�M�{�b���=�C!jo�����Z���1�=;��I�1{%��;*�����钆"4E�\T�=s?6���t�>m3\�sG"2稛� ��~�3�<o�"�ڷH���ܸ�� ڊ�MG5���������������$
�+^�	M��k��Ȥ�3xKnߐ�@1�Ft���{.���W'��B�Vʧ].���Q��j�ԯ�8*��YAn��}m�AG�1I�����Wށ�a�^M>3%%pJ��2�;�B�ǰ4��JjS�b��eѩ��]K"F|6Tq�s���k{�xо���7��?YI�& ��/�'ܐ�2-��ۺ��[	�,{�mݛ�>�`���%��e^;��K��|��e����&33"V����~k��x}9�͵}�m�H*��lHP���ݦ��؍L;�Ħ��[���ޝ0�Z3��S�Dco	����Ġc��DG��u]��J�V��I<����jK�^uM��+(�G�E���K?2��qǸEFK��և	(pp�g�\�R��\�8�80v�]��[��HRp�~�E�������ڲ�C��q�3�GZ����)�秺�y�:C5��"'>8���EM��YM0 V%c���ʭ�����k�����DSE����j�"�va���w<�-��.�>�+���^�>�o�1�k^�����GjG��l��6� �6zQ}#�F�X��}����T�z������"_Dk�CK�v�q�6_����F�F\��s21o�d7�]xڔYP�#���1�՟1D���]Q9�U���c֌⡽8^��9��(����\/��s�����0���a9���Ps����r������U�ZA0��o�ോ�������|�	������q�v:鯸8*]�2��Q3����*=Bp;>Zb���͂NM|����MXn�6,�<�_JK6$��b�d��w'%8��Ob �?��\���}�d���8�A�=�,��T�l� �iۛ���7g�k�˭��o���"+qe�����Q���~y�SH%8��"�]�X���&'#m����B��_�+�\�G-9�0��>�$�9�3u6���k��|u93](�/���;�p<�@�eT]��]�*��?;�g�<-^��I;@�rwr@��M�(��X�[�E�F�SVT]�m�v��]/�$P���D��5J3]{9�5롋�ѾV3��*�J��{=�~�i�B���u�7r vt��_��n�H��O9V��̩�f�݆�Sۣ��ec[�A�!?W��LꋖӄP�z�Auz0/{�9JC�8"b�9�6>ի�3���w\bG��m\K�	�}P��?�t�f�;O�N�F����� x�v�ڥ5�`�Rz����+@K]gJ:����4��&��I�_ A.s�{6&�!&��-�Ȕ��d��i��#͛.�-���&�f�� ��_}a�3h����wE�,�3j�d;)S��|�&W:c�T5���1�̳Z{�š�ʛ��/�"���e��E־K�(��F���J7Jl �ʈKf�t	^��o�B������ �yt/�Z�C���R�Γ�h��نF�ˋ�6�`g>:w��i��o,*���N�*�*`ǰ�Q��` '_���������{���	#CN5�>=�N�ex�\�7j�}�AD�:}ѷ�+�2�%We�7Bqى�RW�]W*M�(φ\��oC��������=wƉc�X+�fbZ�z�b����ȓK���ס�N�Ԁ�uM�˘e�G���l̷?�U�mL�����y�Z�L���-�؏�BV%3�*�ѹ�a����u�0q�0ޟ�<�a���˄�/���@�#2/�8�X�^�p�0)�t���y�yq�`��9dF�R��3�ڟ���	��=�ʀ�AK���6�@�E�9����Aӱ/����l(��ᢙ�d�:�\`>	o�A�U�V$Ҕo���tj����g2���qT�h��:�z'��l�fFd -&�y
R\�8e�?�9
J�]�4����o��W��#r�>L�S������5��0D皼�S�	s�Bk	��Bw6�v`��B��c����s��%����}}��lzp)���b$a��5d�v����Rz��Dv���O�?�3u��Frf6�kFx�l0-�*�'���$���znӇ %�^�ɺ�[(C�o�����i�h��c�{��iזu>���?:�6�z�"g:�p.\���=F������ȉ��"������ƭ��}��;�<��"�)7@(բ�$����@*V��m74ᓅ{=���I��@�����3QC�*)�مU��G�_c%�����1~.�yJ���U�?�͑���wE��-��8-����yR�j.���.������5�UR{�SbG���l��fޜ��ߣo+~n]ٶ���l��qYP��w�;���o�W�x=r��*�%��J@�C�?�𧅶�caj���!֒#����i��-\e~q��Δ���MV-QP��;ϻ_4�Y�-V����A3Ci��Xi�0�E_���|����Y�U�
��@7$�AD��j;�lO$��=�%�?�M.��ɑX
RD����^z�32��J�77?2�8ެ��R�.��PC����֤(q)옘<_f���r����].l���Tg	��x��I)T�K�y�M& ��Q����VBi�x॒ޘ�N�k�/�Q釿�N�C����75������X��](�;���<�Vn�v�?�;�ٝzWәs��������'"Ld�;�Y,�l���ˉd��\�`% U�Br���;�4��`O��#��Yg5H��Zu�"2S�7v`�E��΂�A10`Mj����"uG2����j��{��%v[��j;�g }���?;H�=��0��j7�J��������?\~ɢ(5����r�ٓ��4��<�
V��Rɾ�=����NZ��.2��lh���]N�!�����C:H���$i21s��}4Z}|G�_ܲ�]����?Mg�i�N.��נ{n5@��A����ILu�!�+;8����3ˎ���#�'���A�N�.W�Ճgly��2Ơ;�u��|v�H G��ʥ���,X�1\���2��}��	�$Sx�v�͹ef�8}eզ$p�r- �嶷�����s9�^/�9�N*�����A���x
?�~�f�x�V`n3y����+���ǣ�ڮ/_���F����^�������k�ǩ���;U'�(�{{�D}����n��C���M,�:/J�V!�@�h�i��9OY?��;�����O��'��2�8i����'��+�����L���mU���+q�'Og�8��%v���Qe�8�pK�ᬛ=�m4�����|N	m���ԋB�Fb����*��f�X,������x���8ƙ��u��U�W���f'�JG�:�G�*���F��2u�F���a���芔̬��}\�MnƲ�
�Ik��ݶx��Q�[��d^�|b��;����I;z-���2�ti��sѱ��p����0��6���l��)�A��>:��ѳj�n�fC��6�~vzi��KH<��[of��R�j3j�h��Q�Xčn���L8�ǔ�BaX[��;ϐY
�]�s�BgF��r�<Lnf�p!3�<Q�z2�mJ%{?QJ�Q�k	U+�vs�C����Ǵg��%z��:����M߲�2#�`A�L����$횑/���ma�@?��ɑ����!ɪ�r+9�0jKOUEl��Ą�^|�5�؄
p�;��|�����)V�Pe����[����x���d��O��x��b��N�R���ﲈ���P'G�a���f����	5��V�����+^q�*���tu�� �ϻ/}�ۺ�D�����nNk��1�jp	��Ț$_��i��y�n���zl�D��_1�r�ܲYT��%�e(9K��^ed����x ?w��ӽ�t�^���	�u/6�C�DCܻ6��Xz�q��ڼ����,�đqs�=|$��҈�[��W���W�k�|��t8�+� �)q�E��g\iu3��e�����!���F����7�7?�O��DU�jW ��J?�M��>�
"zHlt'�Can�
_@�4�IA!W#�9�\to�,r�+N���m�����P���'����6U�(C�10��q����%$v�Z�k����?pIv�|�g肃�`�3�q`;�c9e QQ�9n��׍]�89�o�F&ȩ^7��a��,�Dј٠�jP������*s��k�-\:�F��Vz+] [�-k��!�9]��5�||g�=�������ug/��=��`���Dr���m�׳��r�L3A��Y�� NW���T��MP�����Y��K������@�c�j��h�����ч��ϱ�qhel�ոV�J����;�
�,2g���z?���R�m�����d���| �tj�Afr 4iz1й�b|�9��H9
Ci�9X�'�[��"Hrʁ�D)��[���'ֿ�{��EN�s�#�nmy���͐U��G�>����� X�s�)�����>�@�jYf�c��؃B׭��*5�LP{�j� s�	j-��j�Yf/�� J�Y����>�^����V�Qбi��_��C����[��8	 �V��0)��W4gG�|����v�Y5����.�K���4����075�x�yn����M=�{��G�
*�HIa�/Z-"� ���VОY�Ym�LS� ������Qc1:����b_�����N��i�	(�<��J`�Xs���l��+��lk͏;�,�T�u���T �W~�S)Ӵ n{�����y��W���m���A�nṕ&��
�����ʀ����Q��*
W%���5�TRD������(HHw1�PC)"��9��s��{?�?�E�<g��Z{?�9�Q���m�i�3-�/����p!����ᾲ�!��Mԫ��;fq��N�?�1�˙%/���z0�;���д]2}��ήH���8�۳�^[�xWAK����ٟ�:�d��'gC�IX�Oq]��@���P/���~��Cw��<��j@r?}���qI�U0JG�z7*�u�8��a��Q<�I�\�r�3��"��TIG���%`�^Z������f��G��'r�;����~�u�+�O�v��g<"no�P�QC�����P�KLDx��F�W��Z�-w��ɻc�����d8�����v-":���aj4��Z.���?�U:H{]�S���&޶(�����3.�\a3��>���N��$.��a/z6�t5�z�EN�XU��&aY3�tC/}�_�9�+����)F�uW��sU���𹃓�ZanE��	�Z]��y�0���� �=<"%�Zk�����Q���Q=.�h����,��Ŀ��?�:��g?��� 
�-���Z7�H[�C��>���<�2�D���d�
�#/�ӸS��u�W��ˤ�T�q�G��$Ao�z6G\md#B#�6�l&S�T�-Z��A��`V�WD��+�3���[�.�y�X�#�Hl�"��v����"�8�q�"z��jk?��~�.�f�f~P��-�*y8BY����m�E��(?�L�	%��y��%��d���s��]:���CkS �v��c!�����rn����gF��2E�J��5s�g2�!Wk��A8���뗿�'�^���=�8	\��.�|���F�S��u�֍\�����,�UfE���&�a����Y�X)�v����_$h��w�r��� �-�u��{��Е��ɱ!��~Gn]2)�pټ�]b�Йi���q>��Q���UN�	Ug�ɱ�3���nP����}�(r[��9����¶tBx�������H�P�� |�#��h�<9+P�l����(]���M��6<�&���r�R�8+��cĽ���<��q_�"B�@��KMOO�5�+����KX���ݜ����,xG����"xZ?�_�v�����P�1�L��'t�n���G
aM��(O���q��\�����z�6#��������f~�-q����'R�G�w���3�`��0!I��� �����5���~�)��y��ێ	�Z^#�E˸��%�_��k�x�B�̗��C>T�~�rogk6��������ݭ��ǅ��Z�yp��G"[�i��0)�(%�4��ZB�]I�;jz&]�5	���m*�l$���ź��{����і��0�����i��H��?����@Ka;���Z�$��<p�V�<�������>q2 �J��`2�.���N-d��ҥ�t���������.~��uQ6��G�Q~ 7O|���7ż�h�:0$_��]1�t�`��w��_	����Ec����g�3��[*Ą�fb�Ib��O���(�z�qe�B7��1���1���!��D 3�a�������/�Ϸ�O��a��r�N�/waYt2}�¬��(v�	� o�Ϳ�r�Hl~��dQ\\ njA�����2l�0z4�р�y��_P��c����(���,��Wի�c��kss`�2�����K�$y�!^�����|":E�n�>�b��g�>=1:x#ۥ �ـ���x�<IIY�Ŷ��-8�PԻ�ט��.
9��RN }�)ͩ&1��F���uօ��n�����1u�b��q迌~�����h=�u�i=��,���OȢ'�Ѳ�>+��=��Y�x�ey��I�7;Vz�l��t%=����Q���|L-F�%�:~�H,�[��%�K㤃��?=̀O����\�]'}�5�����nzL\m�Q���=�0��Q��-5w1X�b5Y��ʶgpi?C���
z?��I}�g��_�;{� ���w����Sa>�B K�s�oPW�=͊~��CL{g�m��~AC=�}/�f�����np���i�5-4}|Q��pG�g�d�jZs^��ۤS=?��أ�+�mԨ��):L9�~�>:W��_��	$�}�WP܍|`zu��s�%.Vc�Lt~���lH�K���[a��Za������l#�qOJ׏��cdl��6p�
��l6����V=���dE`kq�W�v+���F��ɗ)/��-��W:�ˢ>Ua]}�=��߈����. ����D�G�Z��P�Ѯ���dMv���[=M���3����@��g%���~��Z���{ַq)(Z��
h�#����|��R=�k�J��(���*��d&fR��}������a{�8�5���R�x}�%��˸)��=�×PT�<��?�F7�C���S^B�*ب31%��"�i����Ti��J�c�nw�:�1c�� ����~�	bt�7�M��,���z,�7셁��3c
 )���3�|�������֕S��XG���2���8�:�L' �Vވq���#��8c��ɋ^ױ*Y h#�@�K����c4/\L/`��~~�@*d]'h�V�������@��b�ź��iS�^�N��z��6�̄��I�K�l;�_湀*3[Wvc�b�:%��*Mu����gg�C�T��s�|ڨ�uN��1ʣkG.!�'����}b䌇�\�f��I��sZ�ɧ��U�{$�a�͕�R'����_��nڹ2��~���ie�;�7<� ��!�0��Ԏ�*S��-��!��8n@�>��R�	��gip�+�4���N� �o�3��c�=���{8y�h*���*������e߿�d� ��K@��KF�r2��qE�(���f��J�P��&������#t\Z�}��Q��[�jx	+�AYu}�m
��;�Jd4�S��Y�:�8���>|� 4L:�4�y&V��y7K�A�F���Y��_�q٫����-uI��uLr��=FJC��7�����P�u(��7A��j���Z����м��!V�m^Ȁ� �F�ٳݎ4���~V��Eb3��x+}ǎ�A�=��_�/L�(kӻhxX�p�'��F�1��3<'c*��7�|�1��*�+��;�l�˿�}Ҹ��H�7�Uă���h?�i��gû)ᕅ�\���Yz�ߛ��t�� 7��qp<��VK�]tk�G���A�x�K_nR[,;�y�a��!�� ;��uȭ�S�!��]��ǁN�ue ���9 �ЏM�_�w����~Z�U�F��E�R¼�$�|4]�l�)��hV��cѪ|��O�j��x���Wl��;�o� 3�M��~�:�}���^�����0չ��vs����=�̈́��0f}�*�<q5�[1�-�YFUd@٬���ˆlʌ�Μ���U�^��.ܼ�� ���yȳ����	�y���'�1�}\���V?9�p6wqi}����aw�+_1�j�J֧�n��UU!�����<�ɧ�v����FW@Lf�G<��Ak{9�!�^�� Z&����g�P����<�zk�(o�ӿ��3K���
�����Y�^��Ex�������
��q)Cݞ%_l��X h=,��	�h��5���7 s��!q�l��v�x 5+T\e��c)���J<*��E6���z��\he~�V�X�H7�$y(�����Ou}1�΅x(�*���ڜ�Ax9и�4�����5���O�
q�8�"%�m2�~��'�om�M�ߍv�_}ոg%��o�3U�m}?�Z Z�X��

o�w!��� ���Ei�@A@`�������_9����ˎ�&z��5��)W���G�8G
�r���_��᥁<�:�um�� 5������Φ�y	��)RB�~�����f���ӟ�\xs&^�����1�A߉^����"�N/K웰��2���Ԋ�O�5���y�tqyM�5�S[9�=�N��٭�tm���h���2NK�~�����8��ׯ��.9N�i�#ݥ5+VK�7:�ê�`p}iw:��i����8���B�K=�5����
��}�I`%�C�
��.+洈[u�zJufi 9����j���R�槰Ӷ�|����Kz6�e�"5��X�)��X�zm�1�F7��|V�A�R�NZ��g@�Hf@5`�l�3_E����3S�O�hٱ��}�[���=�4?�UU� �Nf<�mVU��|��������т��J��ZW����Hmb�A��y���)Ν8a<�4�5�Z�iH[ɦ7 @�K��	�����q��!&���w�r^]p�|8����������'��p v�c|������W��6x�_���_M�Y�TN��g��k��RX���$�{v;Тa�u�{pH�G\���U�m��a�ݴҤO�y�׾��s'�䔥B45�Ϛ���<I �J�� U�
��0��x}읏kzdh|`drfƷʶf����½� 3�Xx�
8l�>zY����t�����@��z�3N�A����Y�{nFt��@bFU` SR?�1d���;��Z�!8��p�?̐���5��,��j��7��k=�d�/~��� n�RA�����*�������>`r0�lTQN4��xb��p�� ��z��k/OJ�Q:�Q=>=�v���i8@�K�E7��ی�..a�R�)e[R��B(�1�����)�����bk�\��_����*�+��61t���1�e�%� ��x+C��`t�������y2Ӹ{�R{�'����.1�扰�����I��~$3���2��]��K��s�Bzo4���ח��w�P��|Hb����6v�Hd���#��0���f��|x��'ʫKirc��۷N��e5s ��m7�aI<�'���$�9I�9�ҺW糺�`O�քJ.��~�x6�w���g�����8_Z,��ޢ ��y@�!���v��(.��7�|0ٳ�����t3*@n(�Eg�)ݱ�j{�׷�Ք�śI�e ��h.[��?��A^{|Z2�c-��I#��[Req��t���EP�<����d�>�jF�
�^iz8�,�,Z���NΉ3��ss�D̥�ENW�W�ͽ�~x�!��ؘM���a��䓎uCQ���ğ�H�|�h�K9��ٵ*͖���� �*��ݘ��*��=9�mѯ��[YMD1�a��?����D�7u���ݞ�g	:��)ҳ�d]�˼������\�a(�ߐ���Eb��$:y���ɟ3��dӃ6� �@��?"B�iXu0!��Y��$��l��Ѐ.T�.z�ELK���E����B߶�8��4!�̄��ՐCn�Oݗ�	'�9���r9�wȽ�=��|ݎ�}������
���i����[����j�cyx��-�m��e�I�j������a�
/Wg4j���8��8K!2g`�.-D5-���ժ4�T��5�[�&)��@�>ݎ�ji��m�/t���5G:H=�����pog�7��϶p�&4�H��V_X����s�>�~���I$!��l�YS� 2u�`�����v5~�?}0:��j��d��]�W�u51�w�����쌄�"�b�y<�H�Rey�_�1Q��q�dɓ)�#�3yfx�6#"��r5+t��̱��f.|�o��7�a�O�GRނ���V7|��Y?�u�$����]�g6E)gD�k�̿�u��9Ȣ���ޥ�+^W�f��I6$d�XN�e�B�,��g_P�Ud�{�����w��g��x��j��t(,�Yh����o_���k��mg��.ГB����E���}zF��`��<p��-���I��2iG�����L8��Y�¨ƽ\Y���4���c��qn���p���F���u�_qG�厀Yz����L��8h��MV8JD��1��.���=����Y����>_�����p�Z��wN�'��^�tΧ]�BcH��52-�%	̰z���f�Ftʕ m�ĳGj&�1J��R��g�;-	��p~h臟�?}j� G;��E���=bae>x�\^'PX�@�c����l�ŷZ�gǇ�<��hZ��e�)E�V�<�ϑٯ/�J�|�P��*�����'��ߧ!z�ٳ���R���:��)�o[<��~}�VT���ı�0�0���OIO���'�R����6��V��E����9<Ulx<W�����~T�f�fP��{��X�����%`{Y��\m�X�0��MNw��`A�@#`�f^݊xм=�4�hXʆ�ݔ�S�Ef�������&��ieIK�%�u���K�{��������Op٬�t��:�RaJ��hN�����Y�A˳���~&s�UE��DGOm��E��71���A��R!�r�g?�<OU�*fg�Kʫ��^�1���5�v�V��Bx����l����c��^�P�?���`��o��:M_�0r�l9�*B�Qz���ķ�(P���8����j%�~V%�|��6���zh3��b�ga�I�;�rt.Y�Tw{��q�|C���(�$��Y� _X�A��;|��M��v�u}Tߜ�q!#!�Yd=%�l?���kT.�e�x�I˨�"2���=�]�B�S�N�K7j{~��R�Js��{��������:S��e��iDK�#c)�͞����*7����Q�6�#1�HINFx:,$�9�.���	�j`�gM΀S�YF���u�oxQ~1���[QqA꾜'��=�O��͍k�On k%JNu<���*WK��M��c���.��(�cM������0���^Q-GR�Rv핃}l� �J}�^d�U4�M��A�P�R}�P(�dF�e��.��C�Т�äXV�����Y�L-��Mx�s'��'!Q�t�]E�<{{��GxN�^��BN6Q4�\g��,���1��gg�lrP��=>�,	�<xP�RWǐ�Sq�%yg~������x�y�,*��iD��b8��<�,�(���H�nL�)���蹞��K�̅�BĽ����k&�/��8`Rh��N��gN��ͻR�u�\K=��:R�x��̼<�P��#�^&����>$ �HG`p���/}Y��r���#H]�$ [w!�Y�%#�������0�
 �);����C��1�#�ao�
�~��.2%���n]�\�2h>�Ax{��n��4TU����fL����=;��o[�^b)�VE�	a��������whʹb+��f3�	M�f��$LBu�,yRBL"@�I<7���/Y�/�=en#i�'竉�~D��877�]�M+͖��;�!H��q�:���[{_�U�!��q��!��iE86���?�ʮड़.ʔ��1������!6|��$;<gNV��x[D]�@�fy�I;�����W(�$}ヨ��ȿ5`��+J�r�����qJ��>����\���7��B���L%18�f�%�������l��ɭ ��e:�.�?k;�^_�a�d0�]�5Y>���i_�B�j��IGl�t���v���p�-��Kv�(�j�_ɷ�·!�|Z�/�+�^�HX�L�W+��c�&��Ck�LV�:�Ph�u���@���ډ��T��F�D	8��
���˳J�����>��o{FnǬ�ȩ��*�y���uʓ�*���������~
X��p_�Jڻ�nc3��df��[K�ҰV���G�*�2^��S���cu��b��4�q�����@&U�AwK9��S�<��l�v�7^k�>լ&�j���e��.y}���K�)̎�����z�K����B:t?R"W����T�S�Y��aqB6p�f�u� �E��ܓ`��%�d����������S�i5� %5K��t��{b��꾂�s
z�1�cG9�G�H���u�P:�ILd�^/��+}�&�w�⑴�����76Ny���_�G�D"
���{cA�����)JHe�ښE��E�Nn��4k�7v|(r�~i:
A����͝¸a�E>�U�z�O�)]��f���d�(3C��F�OAu�Hʀl�ա��1�0����!�ooh������VO��rs���d�ʢ���:(��&�'J/�gr�c������Q�*-����H���|<}%$���>��PQC1i�<����*k����[�{	����g�d��1�C��\�*����M���S6�P��b\^���9�>�~�c�̫�G�Ê}�1��W�2��OB���:D��S�=�zt"�$�{w����.7~�H#��O��x�_��kУ�S��ګ��ԓ�&���L� #88 �|��:߿����'�#tdƤ��tb##7���^�9F�ȩ�h��'?A�Á�Y�3� �� m��ϒC�`h��^J�+a,7.7�[�6=���
_�r�1�1��6�a��li>���~kb��͛j�TV�ʹ�i�nl������̥�H�(\�k `�1���/�2ۊ��?�ؕ��=ü�Y�*]I����X�V��<<��o:�=R��ɥ �w��qm:�ž7CD�Go���yS�`]"�Uޚ�}^����5F�R��y�-��}9�`�����M��#;p��\9\��zz\�6���p5/1Lȉ��gNDjB�C�G5E^95�䔁����q��TW��dC�32Gnf0Hʎ�?,"��.��c��44�%���SG��g�'��_;V��*�g�$�>��>��������(U?e"�T�'
M�ì�@�B7�u-�;dVR��?��&�m���>̴�=�yɒc�V�幋phy<�>�����g�+��Q~�K�f�2�l!Ʋ����bl�ni�Rv����>A�:EVh���n��h�[�܍*;�C��h����Ͼ/r����TP�{T^@���I��:`]\��?�P�
eT�G�U�~�����L��~�.��! �TК���w_�S�ʴ�J6%+{��=�Lc���"g��=	��; 2N�O6}�N9Y�I�e?�����AhFG0��9�]dd�ڜ�z��n	�*r�}Cc)����R#��_������KӸ>��4泆����*���PA$Yި��c�@l�YQ9{J����k� z��US�X]*���b�G���cS&�JΟE�Q7�����(��MB��!&TPM$�>U�ďT��R@Q1"��������'Y%Ś�46�0�-�=����� ���ݓ�g#o=���9X7���Nj۸�O�'�(�'����ě���9\�����o�x���j��b���������5��P`� ���Xz����y�k�&ʵ��)'�Ŭa��ù(ޔD��KN�nT�K햋7�U6FY������s��`D�l,��%1`�R'N����|a3��Z�.�v3WkBg�n�V���%2���]AW���]z���Z.���J�����T�zO��H�����m*��%Ge���@�c��<�,�b��P�a���}��q~� �7���-��MdvJ�/b/e��H ��M�?(Φ������Q����Y]�`��k��p���K{>��;��<+��n�E�pu����>"�$�~�r��p/��I�Y}n�R�B�s��j
W;u�z��X��|�/�����O[2��;U�H�p�����a�V͠ AV�S��}��ۓq㮺jI����+PT�:z&�RC`��qL>a����e�Dx�a/W>2~�_��	��ڳʯy��>c��V�O��H��;ߊ��� $C�bo6� $́�j]�Ǭo�[�Sep��|w����MC�LM�EYػJ'���2u�P�c��⧟I��YY�,ڙ�R�B����u��6U!�����w ���E�|�q�59�!95����L�jj���a�	��w�a�Q��D�W����،��H)9��5	�9[��c1���ъ�.��g -��D0Zs��3�Y�����#JŁN����gWD	A�m^�Ī
�o�Gl�w�=}g��b�ղ�ћ��>ɓTd�U�8�?z�c=�&;"v��������|��O  ��Ж��MFe���}��Ϲ5�T��xiR�cI�:b���cb��J�ԸT���'<����9TP�x��q)���D���o� E��(���*�v�/uw��0���t��p��P����Os�2� �k�
 �U�٪��'GR�(�X�:V��3��ʆ�/��i]��ɏEY�hx6���3���Җ��F٣S����ɏ�B����o��˧̤a����z8�8�;�|����� կ�C��cDB)��yr])� QXu�԰E��?j�$:$�6Vݧ�w�ж��������'��@��4��5h0��
<\s�,�"�=�<�%��{@r4���5�N������H�.�ǐIJ ���.�lһ%?�͵��|��f]��Ĩ�K��8[@�Kq�Yl�%�ɂ!8϶���g�:pF�
��
о�Zw���3�N&ԕ�Mt"�a�r�#�0�P+�ME@�}��Ia=�˚���4ݟ�~�u�A��YG�'=I���@%�+Q�h����,�O�&�B�,ε��#����t���)��������~|h�^J�4���.Bx�MR��!���i�o�<�%;�K���q��d��>�T���,�
�jX4���}|+����5OhAb�񈷥.�@���4�G�B�u�-�
[�ξ���e��c%Ph�����)�T����S��홺Ӕ�/������4���c[��}'���Z�f%�l���\����彵���C9�Ȓ��`�x�c����kc��x�v�/�,��k7Yq=yņ��}S�1��t��C��f��^�o��J+��=��}�g~���T+���?�C�S�a��t��r���&^ۇ��Q�4�u�_�w��f�>ʯ��	V��f3|rJ���d���3�R����a�{�e���9{�E�����ܑo[�@�,�="��걺[D��]�Kk�]�Yt���S��糇v?m��{k�[�A�%f����t����рZfa�iyZ{tX��x�(=y_7�^����y��r�� �V�d�Z�.GIAQ�6C�(勯U���^�g���h\�Ҝ��Pg_�l��4F��mɵ�b��%�����i��jy�aQF����AC� x�I�	�A��U�^>�+�W���P�G&64ꂠ��&���]�����&J��j' �Φ�lreg�!�Ks�Md�Z='�CPK �E�N<��:�٦�`���]�nfc�&ﺥ���|�{Ub�4Q�@���j�%/���v�~bk�A���/��]:�S ��e��4}�B�4,�xJ��û}a��k�����;��j�q���K�5�^�Gw7�ݻ�58��g�w�h4�n�(���-���<K�C;�ˋ.u%5��:E�[���Q��S��1��8썵(�V��7��rg��{uKC�����+f3w��Re�k@_�����oj���)vtZP���w�+@n~��E�5Au�E����]�s2:��|� �e����T�>`Є��t!��L��4o��WT Qrm�h�^V���<�6)�M!����j{ud�u0Kf��bW%���\r��� �@�=�|��M������YC;����G?:���VN����
�r��>}6���XNPY �4���˓����(J]THs�zN��{#�_��w���Um#d�X+��-� �:�v�$Iw��\a�0m��!�]���
���%_y����C	��a`kSF�m�/l�8:��!��9����2�I�������]"�?��"�)����"i�j�M����l���]7S�>�� �r��� �*�] ��_���coaܯ܊eiʟ�,1��Yn�c��3�����gL���R�%���,�z��r��0&� .��<Q�~��@k������y �Z�"o�n�C�yqHŏ���uT%@�n�T��v�G�'?�Ss������N�x�D ��� 7�*�Vg�X��jILt��z���׫F"��aJ�S �T*��yz9�WkC�Y���l�{!K��w6��nv�1��U�R��Z�]Uu�]�^X�I��[)��ݾh~�&�!��#@�so���ԕY��g�Ϻ�5R5�1��]E�l�������H��uH�t�5�=��R�rs^���p�h����T���61����i·K�B������n�Q��,�qҗL�dᰔ718��ۛ��n~�K�o�.`��>�QP�j���J	�6H���m��Gk��߆9ǰ����+i}x��i5+W�"gΧ�TL�	�
�gR5��/�K���/�"�5�(Q��'�������R1p���/�rL$3l[*2jv��$rF)5n����|~��|ﵶ4hx������޻���h�L�P��M+� J�����)1T&���5h�8���a�z�QQ��(rp��Ɵ���I�)Of��F�����ĿIU4g��.������<x�l�x>�s�����/Û�f%eo��}f�'/�E��V@������T9�K~2n��<�th�����H}����ܙ/y�b9e��c�H���s�����0Zꡚ�;N�|��^�L�mh�~�\�'`䢋/l{�ʻ�d�>��N�sPpK4*�3ˎ#��j����G���rɢ�lI�[�����N�đ4d�� :�ڢl��u&��r����� �
�X=�4�Wݜ*ѧ}Bhԭ�� �E��W��0��饡�r7i�k-_G����<����n}Z>��B�0��e�o���p��8��p�'3�J��I���V����+N?�;≭K��p�$�h/7�cs�dvp�N�U���Hb(+I�̙� KC��9����h�R���{8��3G�Ym|�.��,��H�Iz��Y��-�V˭!����꾃���k���#Hp0���P}iJu2����j���/��M���u~_ݖ�\�GLt���?�\ǕL��G(����>/?i�#�5#GRG	�.�Tw�<�螿���R�&]X���r|^T_��&{���hS���3@���f���c��O��R�崤I�)��;���F�'�|�SSB���
^p�Q�p��h���S_��D��;��!�;��s�2!�zߡ��l�;�t����ى���T�V6�p��#|�:Yo����m�>)_kB���k�\X�=!����*��,��ߡ^���	t�֢���kRuu�d 9�������R��w<��o�[j�F�c�����1�P�U릫��`n�<�t"ST��1��`Q���6�L~�R~y*�%����P���&���5�X:�Z�Vqkw��"�S�*�P�{K�!#0�����	���A8����;U泆k��s��)����%`���������oũ������q��ђ�s{rK�F7M�0I�n��vn�4�^���?�ׁl@tFe��+�Ŋ��T��*��>�%�+��n_mn��p��L��ס^u���g�~�-7^Lp�VD|��fM��£��2Ax]�n�e3≜ܲ^��������Rۡ�zzc��v	�;8�w$�&�zɹ�#}<m+H�l%�q����Q�I�����$I�8:pl���>b���ikq@y?�t�Ω�h�i��-�`Һn�d'
#tݩ��fc���HrM�=�1b�l�J��O׻49+�7ŭ��9_�q�&�C�o��+�*YK03�Np�bG.���&\��t+�y��7ۋ�"���PPP�p�����P�._�fc���tݲ�Z0�NK +�բ�����h�(�ԛ�Y�d)VF�hMY���1B�	N&#%mM���(%z^� �`��R+��x���ᄎ����Z��v2�C4�>qs��?�!�~#��ϳm�R�ڰ��/�Wl��V�����9L.p�=(!3�(1d5��6,�>��%�������L9.�o��Fp��s��RdG�$���R�A�d� ۠io����x�\�e�����$��`�ɑ�Z��q��vX$��/ܽ^S���HZ�r�M7{|�>�?$���g��z{��U�a����Ma�5J�yM#/{T�|X5vX�8s�l9׾��F����3���!������|�5��pz��2��˻���G��L���!@� �E���d]�j
F�i\˽Tx�@z?y"#�P'�V�Dr�A�"����ZZK��	��P�Oh�̡�6����s��{�r3��]�㧷��uG�Y��WK�\�C�p��6��)Gb���`w_��)��~`S�D�z�m�l��,�}.�Z?Xqpi�%>2L��6_� ��+KV,#K������o���7�˯Ҫ���n{!����H�ҜU}Bܐ���G�q��],>��F��e������n@��/'��Եg�~4�
������䊥�`�V�u7��
���QF|	?�Ûl���h�����/v�1���ox�6N�<Q��P�s#j�l�|�ܰ)˘�O"Vs�We�f ���Sf�շ�h�r�a�Ks@�3���2�X/#�ܞs==4j��y�4)qimq����	t�w���������p���n7�}��4����=�ᒊ�5	��4�RXZ���h�ެSh6��fʅ�C���;��[t~�Ī.�}���[�AB�JƓ�vG���=�P��F"avq�b��;�u���\"�Y��d���$�l�}sXK:��>Z �bT_b�:窇�F��p��H�?]�_ۋ�}�����G͞nJVX]�Q�/�Zfe�|Z��������+%�M��w�݅�}� B�C�Ն�}	�4=S��r]��C����$��������q��J{�Yb�������Tl�q��\�$V��u����\}5�+�K���uh��+��(U��B�R��Wj-��(�ä@�\FL. 8�vY~��������^����aA8kWH=���� ��t�y����W]?�0.�4]���1�U��Y��
1q���5�g� ����%�Ҹ��8�q�:�����*��^(,_-����p^b�P�e�/C��t���b&��V�kڢ��?��!��L777�iJiq�\���	DV����w�W3��� ﰑa��O,{�I���I�*@O0�~���I��#�7>����Tͨ�h��d��vi�����+���N�֍�%� _��ˠ�Q }S;D^��^)=y��!�%MY�[��Q�Y�)��=�cE�g-��+H\�{.�v�_��˓PZpZ���z����]{�1�����LI�-���]#�fYJ�t�����{[����VM�!@��|�mu�uf>�:Fɏ���ZoZ��+O<�B���E3w	>�1�v�	[	�����K�1����pz��wmyT�F�m�{;B�өׂ'�d-?������i��C�w�i��V�	��N�T�;�$H
J$��cP��3%ˬo�f�\�?]MqyA
���s��-�#��hC0�|KWy����(��#-�Y�� w���)��Q��P�����,��QP���	���YT�,�`���p��;=��?�J�EQu1�
2�E2��Z�2�ֹjR�W]Wm���A3�QZ!�\q/�a�>�HE�2uuX6g�Q���ִ�4r�]PՏ�G�p�qH��4��{?K�� ��T��TQ ����#\z4ׅp�<�Ѡ�����̠$�wV��cy�f�g[����"*I���(�(�>�aj|�gؠ*C���P�,u��_!�^��T�U�͟��?�+&&Z�䚳^9O~����<���`��5y�B_ -<���૨�E^�v�7-%����p��5�,��x�,m�?��	��;��G_b�����ʳ6����4���۽9�%��iCq�,Ν�x�G���$4�Uڸ]D]0ݢ�%z�e#FQR�-��nm��>5Q�rjq"�(�d�P3��ld^~�d#�1�:�9R�c�<.;vjjF��6�{�R�I��aɔE[��8'VBn�
��k�����a�U�#ul�����u��,߰e�M,�����UvO��"×tCk� ���¬��"�;��!K"���:�	c���W�Ĵ�-�:%�HW۽G�0)�����,'�-Rqx	h~
0���I%����k�{8�y]��e��r孲B��K����>/HYZ��DS
C �&�)z�N��l�Zih#�ޏ�U$� ^cmj���TN�'��w T�.y���d괹k<���SSĔ>��L�I�La�I%am4��ު��6�PA�f��K�u�>���pEG���Ϡ�{��H��KI ]�w��;Ǔ��~!���.�lo�3\O�Ͽ3�x*0�������K'�fH��D��	Y�r�S�f��� X�D��:n2W~����=�uBڮz�8x "�V�%G����+K�@�e�x���ͫI��7-H��'�]P0�,���@EkY����7�?��,��0�Qr�����2@7m���n�B����zVm�T)��dQ�M').�k\���;\'��n�[e�fa����,2<A�,uӦY��X!n(o�Pxw߽o#1�����A"P��u�InL\���.�6����ʜ���o?\؅E�
[K�a�'3�������v�289���Y#�����'fI�(C�<����T�#���rԜ"�8 k�����%n���{ޣ��{`�ϱ�]	n��˨c�:ol�2*g���y��}֨=h{֌�"�6w&���2��w>��H���$�k�����c?#��>�����}p���j���找v��-��)�y��-B�QZ��{�X�V�&_��� Y�Y�C��?âx(]mXFr���/{�.R��B)aH�b��rV]�����kT��3��D���[��MU�b��ŉ6�ʱ�|���٧6��׵�����lU��j�a��<<9H޹��ړ��[]��k�K/?�g�W?� �9��<��Rv��u�+k�o�Lx.�X>6��w�5�g9��a%�U2�4�s1�},dZ��:M����&J�E��zlӮbI����7�G�ֳ���7۶�@'ݯ��Ul�?;�ݓ�hl4�"�h~ʝ�4j�q�(Z�q��yXPN���&�!p�}�U���X��ٜ���[�)�/�ӿ���[�ve��������v~^r��C0"I�K�t>�9�����U���i�l�HJ�M�P�����I���dC��zT��@�8@:̭J}���X�c�"չ���o_:7�0"��h�qѶ�:�1f^w�R�i����(!�1:s�5�j��h�)�g��x�c�e��I���Ŏ����h�#Kp�G[ 4��c͡4v!�.:��
����ќ�r�aOs��R1����X�k����\F���v�W��Qr���Ob˷SN��Ngʈf��^��������C߶0a^u1 �6@�;�Y���βJ1�6���5�u���jKCc�	��2�M� ��|���X���(n�s0���0�gi��qE�������t~{z�X�N���U�{�k C�H���4o��Uu�mq�NP��f)p�OdXs�@����E��Η6�F��CK)��*Fџ������=���/ZB��DO��A����}"�{e�	���0D�����=��;3����߻�͚���֜����g?�{�3�[��8@�Ѹ��N�����\;󈈂,��n�}ZA�L}G����:� �~�/`���Wө6�h4�z��Y�K�p!��7�SE�����P����B�٦c0��R�]����D<����j�9O�J��a�蝥8>�iG�t���k��"Ü���ln����AC��M��kdG��L��+��������M'�i�Ñ܊*�OR��i�64���	�.�;q1|͖SV��gM
�ufKi�E)�����\�|ٗ��C��!���My�o��)-_%���w2��N�)r�Q����n�!�I�5v)��O��ۓ%���|췮�ܺ�4R�bm(]�%�ta1;���� �;�{~F�1�v���*���P���g'k���9jAK��jr��l�;�eN[�E�9��9&���x��T�[EiN����РG��b�Hs��-���1�Al�:���Or��L����V�o�l~fx�ὄ�e��UG�����������P��Y�7�������}n����p�����Y5h�?�u.&Ӓ�b,x��A��`��E\&��)ZO�y�_w
6�i�<�� �J,F�9U@Ǚ��A;q�x�j��u���L���3���C)Q�>����=ظ�vE0��ei5�VA2�9b�5a�b��L��
%��A'R&��}iM�h��z@�e��@��@�[�,��#KV;Dd�%+��Ľ�z����t� W�uuUi�y�C=Ck:����sj�vd:-�{4���t�7�p��S�2�R���szM�'0�~��h�j�$�U��&�hA,&��7�,;T /Eq�O�`��k[y���0%`�2�gf���[�_y������w�����v0�\+������ۺ���<̃֠���	Ʃ�U3���Pv�w�Qd�&�E�q���� �Z�� ��"b��L4��@t<��&,���# �ܡ�o�5X���Au�2�-�b�?��P�����¦�W��1�pxXb��ޣ��-�`�BteX�oZQ��Q�87;;G�i*�~���w�ab���b��}���C(`�ؼϕa;iO�O����s!�,J�`c����m�B���Y�� +��?�a�K�Q(Ts���(�����֪m�қ`3A�ȯN�Ϟt�̩Ҧ�&����P]:��X�w�2/ �`��?.d{oH����Q_�Ť���b��q��8m���b�a~�g�3�Je)�
�,��`&�@+�NB�%e}�bu>����_�]|�0-1��K������K#��$�!s�kk��؝���뎏H�/UVZSO�`+�u�n��h�;�-�^�}#6�Lg!_z��^QB��5*!���[&�:f�e�]�%�a�m��.E��C�����|��x��@�DJ�3Gh�}�^�GL�S���WJ��\�[)�<v���&���U���;8`u{մ���c
ω1��6��אs�l����˧B��
xTM���SQ����KS��	�PJay��>�ߟ���q��L4��U�E�\� ��.� ��jqJCy%�c���"mfj�~9��%^w��#�q#�a⹻�.! ���|>�T�U!��mI@Z��Q�|���IB�~o$Z����uQ�ޗ�Fו�MfqsY4���Р�c5�Dw���O*�	E?nb�k���[�{ٗ��7��{��tuU�՘'�ߢ9}��A=�=��Յ;�,"���N�z�@0���λR�u�$����5��h�1{.���Z#��5ź�j���V��z���d�d��++'�,��K9c`�?_��]n俌��Ւ�L�ƝƸ�gu���}c��r*q���f��k�e�u�@[� ��!��S��!՚�T�wT
|�*�;Wx&�.cb�1J�k�>y����f�N��~]ʤ�&�z��հ��P<��i K=�W��{v�{�_5g(9�&�6��a?�˗��|?�kɣ�v��jbQ=�L	��2���׽J�]6a���.��E�v��CP��-��J�v_>�ݢIh����1��0��Ԯ�K���EJ���T��(כg�'4��۝��_���m�"�V��мʆ=f��+��e�ຼ�R���F��"5�K��2�2r}�͸�G��y��E1�S9��˘�T���jR��z�e4�2;G�N]�3'99'���?��gSf����� '���h6�{��t�ϺD�	RIO�i@���CS%.|�M����bL�s|�w����!����s�K�h�I��l��K�}E��H71V>̕��u������E~�(2� 'ac���j�(>�H5���1���OJ�����+�º_^�1��%9���@%;}A>�-7�@ �Z��?3�p�SI��.�n��:Ԕ��*u��H���+O._�<Qo�&�i�����K���>-D��Nr�`�'�V��>ޑ�#��7˖��b���s�ð�����<z%��CΙu'��,yV�b!x,e��+���Vo,�ǳ~Y,K���@��*}�g�( �ȷ*�:�\_��5�>����٦�p��;�[��U<�n3cתE�C��
�ēr%Hn[ոN�/�|�s����E����H��C�USM�lI§%z:_gQB��|B���b)��p������X�[{���3�3Q�U҄���o}�%X�I�L�^�@�l���w�a"#����sU^3����a`;R0!��ٶ�2��+%�5B6�w¬N�4�;<҇���þ�s��-T�+��t����,�%N)�E�O���<�
�ؒd���6�̽��ᶽ��rn�!��:]���W�}�p��6j	5��&��� Bs_�����̃�ً�����|����&쎏�ܼV|z=�>�n^�@:s���mx"���=��U�F�������*�^�,�d��Tȧ�p6sHC�ښ�J�j��c��P��_H7n��Mo�ؐ��m��<�N0�-���()����o�[4HI��Ǌ��L��=Wj�[<|�����	��K� 
�ֽg���æ�tE�R��|������\�o�7�7���}�läRP�0Ffa`*��aǷ<'�H�$��D���}^��@T��Ka�{��t�kBK9���+���`j��JRtm*�<�y��Z��d��uJP0�f�ペ�Ⴍ��L�o)�b��Ht�w3���#x]������dj��԰7lP�&�۞�^�Uu5��}�Q��gi����C��,�V����~�`���xv��;%(q�����Z*���'��:�Mps:wz���	ww��3�kXb��櫎21bJ�w��]&�"��I��VYx�/Kè:v�߾/w��V]��(����뉣o߸\)���*��=�Fɟ�L���.Mؤ���N�Y*����\0��l��P�a�Ob=A��چA��A�<�?ͻ���fU�5_0˷�Ȭ\d��m;(w��|ifc��R3���a�4���4I�K.�Ʌ��݄O�%���q�~� �v�~��ܟL��|�ǜx_����y���L�m��_
By��btN�=¯���� d*��V\5m�n��mS9,)�%�y�alXm2��G0�A�A��b�<ޝ�(��3�/~��� ���J���/`�������uO�T�%*:�E��f��bGEOD����*�B"��7��r�J���\�7P����t�Yk8\W=��ܾ�+����l�r��m�*��ꚟg&>�9�����%&5Iw���RV��b��3z&9X^&t{m2�K$��o���m���ec����r����cD D�����C/���5H��*W4�,!�S�!�Y8yP]}��QV��!�U���%$�w�R���0��-9�$8���)ǰ�����f�ꍹ$�H�����a+��zҫ�s_3J�?�B��==��QJno@K���3��q��̃A��GG�V�j_��;���I�F	l�r�G�М�3���I�Xw ^G��yQvqE�M ��>��T�G���ݕ~;�����Z�Z�^�����'�J��1S�k���Q�Yu�|_иp��d7' H�WT�ڹ��﫪�F��5�d�������6¢��ӵ����<p�\W��|&�5�T*N�v[�b�V\_���O��h�l�O8ܶ- �%t,Zt	�[X+���v�����\?�= �u�(�T������S�4-��~�+^ա��~�����ctO�ſ��lc�z���JJ�L��kEO.v�����#<���u��$���ݚ����O��G�ie_���?�5�|�*��.�{d�[�O0��b���;5H�WH�	1��w�]�'�l�ȷW���kI�0���'�>2Qd�y�����ǒY��y���rD*��<~v�� ����Cd�#ث�f&rb�Y0?�hL�ި�����<f�����?,%n�����ߵ&��-�iAz-M"1%�x��8DV� �m�nJ�F�á����o������N8��f�]�Mk7_R/z��Z{��͕Fx�������b&r��+��U��ǽ�z�ܥ-�'u܉��Vs	˿�MƬ�&�pYl%G1���cJ���L��	����l����W�sR���D������N9J��㬹� ���)��z��=n	r�t6�&|�=�.��n� �ͬw���Z��*�uz�j�"qK�v���M�h��@X�ǽ�׵�o�TV�szZ]R)W�8��,��TWy<��;e8Uz��W':��!�P��0�hgۇ�*R�EI��F�/n��̖Z����K�N0���ğ}�ma��R��at5~$y�7��s��Eq���4��_����.OE�<��8E��YJ�nȣ\�D57�k�W|�h����P��=�J��PV���:Keh�T��6�TS�7 �����/���פ��*��rfPi�L��l��{�^\�	c�2mour�Ѱ���M]I�3B�ϋ&�!?��h#�&!c��e*��OgD�4^�J�����������$�jW��$p�љ�%���ü3�n-��]�mq�IRLUQ�N�<8q�#�̈́���_��_���<~��M
��l��_�C(���7�>�V�0��*?�׷g%re���6������ߍ��3�"��B� }�Hb�����a��Ǒ��z�������EY���&��`��ٖ���}̊:-�LƫyH�`��{C�l�_�׽��e�8�G(�0jSsBto���jk�	D!��=���]��7X���z��9���f?�fw�ɯ�-��B��tƐ���v�ߨ�;��ڪ��IB-�*�I"��AJ�&�r��6������oJ�ZL#�[~�C�/�̕{r{�<�/�|U*���\��'��������j=�@_�����0����ܰ�e.BC
?����H��4i��M��S��X�f�82���̺�6q���>]�v�$�-����X�]�U^�����|��d�z�I�|�}�Uw�����W&	�X�%�w���#6QlˊK�t�[Kƻr�����u��Ԉ�m��F��kZ��t ��E�ʐ_�A�a�AA�7���Ӹ4����~ޑF����a������#7��aߔ�x��z������(�-�tl�7���`���,�b��P���F1慭�b,5�ݳ�>��O�7FڏWV�S���\ZXX�0�#��"*��~��ƙ|��x+���,\Æ�c�K�Z��&׸�jX�]����� �_MԟM2�_��#�u��Xث�ǆK,
�����wO�HmH|���Jw��rf�����oe�}��Ȭ(���xJ�hM�����$J"��aч8�<\�Sؽ��.�9nl1X���@df��o&.���l���{��Pq�6�2����Gx
���n��&�����1(J�0���1Qlu���l:�e(��ak)*���&Q���#_ӁEǂV�?�\��Э��
��9Y�~=�p�l���q^]��~�az������dvT?��,x/!���/��<��1UUcee�v^$*�[��X����j]Xۉ#~-%תJ��I79�պ��Z=�.!�w���K3�Xy���y� ���/��un�Y\���&���X�Y�4E�����cu8�-{�`S9�������Z6S9�����3��S.U}���݉y�	z�^��k�`)��8�
>�ޚ�?��m��~��������@A�k�<�U�5+�1�*�=#D�}���!�,�8�s|�i�D��VC��j�ԞUt����݌����`�^��s�� YOY`;K�pФ�CN&@sAt�%@�5� �;~��DZ�iI;�����Ӻe���g��{�N�S�[^��x�d.��LDkY���M�\��>�������qN���&8>X����V���T@$�٪Ȃ��O�7KJK��Y������
����������1��\�����h���Fգ�v�[S|�J���j�U�����Enf�G@i�d��ԃ�ݽ(��J�^pF9>�L�>�2�eJ�=�<���ka�]�J;l�dK�R�\�Yb!�a� ?Ĺ/__����UӜ<y''ϣ��(v��j�є����^�O� � �)�ég̚��g��Q)_/�m��y�]u�mT�A�ˡ�	bQ�����u{yޞN�|�mS�d���꾋SP|H�0AJ6<̴��Q4'gpP���nj��mL���I�`�=Ɛ�ͣŖvR��"��`Z�n�M�v��od\�fS��0>��<�I'<�����I��� ����#��<(�~=����w[Z蒰���ܳ�a_��9��]ɞ���wr���b���^J�,���l}��z��:1�i+��t9��qdq�5L5��/*rk�ЗdhV���(�d�@�H4XLV��lQZgs
bE����>�}�=�����-��ѿ�F��6 ]�'����?���Nv���~W�tz��֛�}ˋ����'Y6���o�Ȁ�fS����?����s����8��r�غBi���q�B@��@���\�;�n,Ɏr\���W��K7}����,�~���Z˛\m%����g��,�Cwsu����^Y�����9�8pc�N}��żN�-[�r�����L�BE�;y���"�
PX���B$������Q.��6�6��+�zi��.�+˙3�g�+��Y{F�/0�� �Z��"GLt�����_����ln�O�Ξy֯+O%���}��[�>%AQ�����ٱ2��L���MI
pYC�sȻ���Δ�S�m�[O� ;j�bD}����6-_|����`�Jû�ire�
�X�z�eQN�`��c/���=X�)�9��Z#�֤A�����o
���zs+�e���D;�0�t.������'3�49K���+t�Ţt`%�Q���ZO~P �f��k��R
u�u�M�W�i./f��4�+�"5CY>��DۉM�B����4g��G����m &�QVX5$~�~|�ָ�X�y�N�)�L�ԂF���̨��n8g�o��U����1�҆l���<���E�m^8O�^��m�i}#n�ڛ���Z1ڬ�9��:�4B�b�r8�֐�7�ˡGv�sT�-(�U���(l���\�
�'I�UɬoO*��ҭ��q��gU��M�b]v�Ӟ[p~�b�@�r� �C�QK�j��X�4q�Dj�R��6�*%2�$H-�/��*�F�����+d�_�fS���dy`%����O�wY�X�ų��9N]�UYI'.�zeE�����ӱWڅ���p6�G ��L@���w�]Y��o�r�(\?f�.t�eq�2�]'K��[������s��%�_~�Q��<�R��nU+�74!�em��Cp�ⅰw���j)}��/ňy���TI�>	��]y��?�(�E�$�pK��ؑ\n�I����[bEyW4��,�z{
'b�Z�╔��z�;5�JԙMN��6�J �ejV>o��&���#]@q���r��6�I���_J��H�{���b���PӍ��W��*�Ӯ	1�4mVz�e��ë�o� i2m��,ߡY���x s�kD���]︪�`���W���*�^�-��0�F�N�CV���_E�!~�m�U.�3��^exU�nA䟸a�C��Qt$em�}�c�V���N�SG�Keeb�K��n��ʩd��핗y�,�O+G:^�G��$Q��s����Nǉ�U�)���(��#1���*��H s5!�=}�{C� Z�Z�R�<d6� m�J h�A���՗�T���:nؿ!L�w��>�-2����d�.î'+���A;M�o�C�'��*�|��m:����a��S��,���IC�����xNR̔]R�n��aE�� +��|�!!u\�wv���2���b����Yv:��/���u/�#v���;S�T���̇�<[�?/[Z�v��@	�����k.�m
�N[j>�d!F�P���`�aܠ���W1^�H�>&�{5�1C�p);E������g Y�\&�r~F���x�}�Kc]ڢ~J�N�X<���Qs��g{�/����TGg����}ӡ7~؟�a����F���M���DK�:W}�v��kpM[�w[�Y��B�&�7����V��)#{�\�����%Lg�$��d����	)gZ��+O.���N�� �訽��\>5�Z>��RG�RYpN�@����mv���k��Hbc��Δ$����(��7�X�P$�����fzs��U���z��CW�ݵ�f�Q��~ܦLE�TV������oUcl'ΧnWk:��$�eq�����5���ɴ��T��:�䊺�s���3ފk&�F"~�{�{����V��>|���1j)��7fP\=���Y]!������y>����~���I����b��=:�s���9�2���A:�ؓ��W�l��wܭ�]�S�i��}��.՞��Q�+������3j�&��Q�N�_E�̟)ڄ��ǫ�{����m�.ͭ���D�]���DE0��"�N�I���L�Y�<b��!��¯�S��y0���'��L��ލ���^�Ma}���5'�j��M�����kw��~����I�M���qg?a���Q��4��|'Lzwn�`�{��|��<;ۀ؉y��C���(��w����YxL�Z|Ǫ������òjֆ�"�ۯ�ϖ;��P��C<s�����uu&ԕ|�6�πƲ��q��P�����y��P��w�e7���`5Jes^�;���m2�T��j;;������b^����I�^�ގ������H,��/z��,3��I�%$?�+K(�~���{3=	@P��ю�� �w[�_��o �s�u>��DM���U��<3j�!t�g���d��29���YG޾�/�=����ek�6h/!����RpNN%��������5N�]m#H1��:�sD!&N��.��pc�?��^R��äH�S�!u��ABϦF芠w�����ɝ�L�o9�}e��9��iP~�x����7��wx�9�9@4��]��5�\Oh�'A*P"����h�c��)q�aH�y钲�Wl����})�[=��zMq��VJ*m�Ϲ�]t|PZUf���.�?ҥ�wb?�&����e���9/~~�faHLAge?�S�
hKZ����^9�":�)e��D@�vr�d�g��Q<L���p�>%����ø��v."��=��A�",̍0��uM¡i�UC�cɔ�~�ܤ������a�֏���W'�൷(c	�G7H2�B����S��Ki&l�}iwD=;栟Q��1���`8]5u�ޤYd1(\�T?�F�ȓRЈv�r�tS����O���1�X�1[y�5������}����5)���+;���Zk1n��)tN"�l�v����m�̧aʵ�[9r������;�ߞqr-��R6{G+Zq��ɢ�$�����\<֟��P��PK��:�kC���&}O�E ��=�[yQc�h��ǆ�]������C�n�O0��qR�����8们�3��Q��j�d�M�Rd𾦲���%>�0��E���]��y�<X�oc���n� >�9𥘱>Q��%���f�����`�O���������b	UJb��jd�VI�4)@�?���0xMo�ۙ%�~��x�
�0�ݲ��-_�\�<������y��J-��AQ5V6�Fs��-�d�U�e! ��x_��U�+"!y�t����$:J����K*���O�u�f�edul�%���o�z���C~C�L�~E"S�����cz�����	�E�/���	z�9_��c,rm-�	��lԘd�	|I��2�IĭǹNb�/.-)�H�ke�����!��b2���`��0{���`y�
�����NDx��s�-��XVƧϷ\8N��p���cNX����L�}sE�I���WlN�8�z�\`�����?��
G���G�ޝ'g�^����.g����|d�z8����}�V���<Y|�����<c���X��bo�$���hT�\���2��M��	y�^��V���O�w���Y",n��ts�U�A�n���m���dF�
��ۥ�.��	�mz��2��/��m,R��_<�m��K��9T�I�ٜ:�������S�-qR��������L�����3(0����P����;mN���U��G��j�o�bz�	�P_I���/�<�}���� X�E�o���楕ɝ�l�23��,f�~�'��<^����:r��G�]�u�2�k�6 �?̬WOl��K1�ђan�[c!�0,�� �J��	�c���T�B_l�]b:PZ��Aa�,;(���7��6��I�7��;<2��`:�:��#�$*����柝�0���ݮ���1��2��B���}&�m������GX�@' �V���gYMر�Vg������=mTe-�8Y�@$��w�w� ���W��I�\[]�=n[��y5)�K����5TrӘLXmWCU(�z���{~���b����?��n{F��b�/u�K��M?�T�7��ݓ3��<#TP]Qj� C����	��m�vCj\�©�F��{&���I�Fq�|��N���Ft�+�̙F����*+̦�i�Dt ��βNg	��u�N`V�_,>S��Q�:ߨ��)�SN���j�Kkf����%���زm���,��|�α\�@���`'���DJESr/��㬸�"e�|�'�����],�[*V!����ͦ�9���Kg��Su�3��F�3�!�-A�bG������O �4�o��� pPw��
�<J� ~|�ۑ�¦$���^���c��FX���T�Dd�U�����)M�"z��C�-��J��:&�0�F�������z�����<���Z��(>W�f�����$
6g2�y��4D���W�q߸�'�Z?t%Օ�"��� �s���2#(��&~B��ͻ�t�Xz�6�8u�����7G��OT���!�.�O��;��G��_0h��-�5��=�n��<�ӦB^��R�Xq�X#�C������@��@;�w5p�K��\p:���ixzy%K��~���=k�6�%�6�ib�~��T�����X��˗�ﾸ�򞎺`��~!Л���Et0n$��AL�G6��IƊ!f�G��?w#��Y>M�?�cӝ?\���ʩ+�M�,@���Y��J�{�m��1�C"e�r\��Og(��96�к�Jo�lŤD�9�H� ׆)7V��w]s�Rr#��n۩꟯�'��8��H�]�Z;
-���ҏ��a�r������������;����GYb�&gG$O��G#�g���$ ��ba����n��cO�/�k�<�mX�	yq�=��T��ә�}��������c�F2�K����bcm-�u�eA-���xD�p�|�-<}w�FU�a"@���4(�^��q*N[u�$�����J$F٥X��=����M�:8x>ZQE����Ǩ),lc�?u�����H拰�N*�a�t�s�t�c]/�2�t�}���88!�����O�	�c��TNn?E�<�`h�4�Yv��m^���h^�iL���a�XlH*���Ӿ�_�������蒝���u��+�j���Ot��O�C�Uc����`mG��w���'N���}�Α�|�R�t�N�Tj7"�7�m�+o5H^`�~H#,B��-���>��7��-1����6=��}Qg�J���]#�s��;�ִ��L�H���SQ'G�V�U� ��>�6����p�l	����X<�B8��7�H�8��h���
4�f�3�m���j��fڔY�c���6�V�e�'ǯ@N��W�7L�cA�O� S���`�)>�)��u��$��Q���C��|7�#�Ϭ�E d������nX�h���q��v���B�3��E�O��u�ylݧ�������S|��e,TZ�zPN,��lw{n˷��Pf&rf���nS��\+��--`���O �=ʎ��6r�0��B^���bb$��7|z���-�3�5��"��H���[ۗ���l���KQ�b��g���<{��y�Q��w^aUA^�׀���u@=e.s��>�o�q|Jr'��re�����B	�^#v��q����Db�K;�J�G�CLI_Xh����b1  hFw���%�dBb�\+��o���f�jQbn>�ޛ�����t@
�����.�g�;{N+�B�݄�lh$�?\��Q��VuAq���N�x[d>�ز�v�%up��������ˤ�.ͅ���ls]�4�mƛ?/��k%�E��T��f��yK� �?������0n\�n��r��!��(���yR����7�Ĉg~���a2����s�5먑�j�̧$-�?�]i��/���eQ�30�.����f�����麼�d�g"�ϲ����M�~{Wb
=t>P|��5� �̎7�ۯ�n0�m��;�+�[& �y`?�:ۻ@S�J��M@�gx{,�9چ�u��k�om��	�)��C ��e��Ϩ�,��҇���#.3��@,U��|@oNf[�TR��f��P>���~.��< lΞQ|�놋�M�,TvJ�Q���H���`�V����mg��"|i�ǃ�4��� }���x�`�gKZ3���f}��?�,s�㵋~��G��u�{d�no�&�wL.q��Rxp��@�%����t����t��2��ϓ#'��4�M.xŴ:�Z�]������]5��x�*���'do���v=��
��q�q�5(��m\/'�&;LB�HM��T`���󜏇w !<J�%���_�/�m���e�l�m�W��6_�x1I	��[�ls��F�e��*��0���?�8��wM� ��5CO~�4�_����P���:�J�����5�0�h-n��W&�>v#CȒFRT���FJV��:Τ 3Z�}�~�7�3�ܡcu���	G��&F��<7��jþ�d��	���!@�:�)İ�r�_��~�ָ��_�r�uw �F�u#ٜ,�(n��|�7I�xv�ʼoe�7���/��w�7{?�� se�9��0Sg6���`�pA�(������G��r���`�M."�g~�w��?�j�H���4�ۼm�J���L2F�"U!��]I�Q��5qj>/�$��9b�!���t|��,����@�Kj*H�4�j�\(����ܖ,q̠:?iN��V����e5��xh�������ve�N��S��߯6��f"�=(S���ӓL��z���3��<<Z��{�s�O5�7k����Y��J��[K�� �oJFL~涹rZ)�a�BL�ۖ/ct��)p֓p+gh�Iw`��+t�<�j�q��A��^���+�|J�;ĹO��M���%�VS��\;W0#:M���}�BF�Á0�
c����;6Co4M�� m/��F�#����:��<�5��KXl8�fb�Tj�4q��m�!�f8M���G��mJ��c|�'_H`�_�/'�OtAΦ6���}燥�����_}{����N.��.h>*�kI§eup���<��+�,�b�.�&~�z���o�>[%nu0���q&ƺ�GQ\^�l���k��N꿋`����,8�cOL>5���������������=��~R�.�Sѕ!��Q�Z��w�r�͟�T��K A%Di�v�ȸ����P�4O�e�)�Um�������A7e7���Z��Q�x���w�4������ן�L�cS��67��/�
o&��=�P��X�'*}���Ϩ���n�ʔЇ�	�v[�q����
cw�{1V"�Z'����=��U+��v*s�Eu,��`u��D��>��-����-<OQA�R���>�w���n$:�k[[��D����{�|
����ǅ^���`~��u�GU���(=�M�d�"����J�o�(e�v��y�6�G
�N�Iz��;�v=��~j��������et)1�,eI�<B�*ԁx`�3
F��PQ��#p�"b��_��Q��Bל���|i_�'d�E����:%��'|2�f�{�u��ӎ�t�1��J����s�5�����l��"�)C�K�5��'˪���M�s��to�D,���s��r?�!&���M��ڕ�_�>5�=�G�.���	�\��'�%L��o�`R���F�q��r�%�QI��7Jk�D���&�w���B���I��i�Jt�>P �mA���f]��^W���o=S��Sǧ3S������J�e��}�ނ�_���; (�M`M���?��?�,:p#j�Ika��Uu�{�� �`�G�xa��b���E*fJ� ��1>kZL�i8��Dr�5�2���;�6��&q'&��u���[�Y�;}�I~�GT�By=%1�����q���wO
]v�e����t8��x�H�^��F/�=9�&��~.|��͆�4�x����Q��4�p*y���(5�6S+Rx9�Yg��*fKp�m�=�����`�jquK�1P����şg����sE�)@'�h,���I_h��p��{3��	��{�"��n���6d�&r�k٭v=��X>D=V^b`��?�ƿ����(�"�ֺO���~��� �,�N2?O+�˓J�bL5$�r�|�}�#����=X_~S��̜ Mb�P�q]���]s�]�u7��������.�S����UP'
;�h"�M&{��}��Q�R�Ƀ�:l�� 
{^gC\-�n�}�F��Ӂ'3S�A�v�D�k���Ɨ�Nf�O�z=�1S-�X]��g���ӝB�`m6�6�C��S�}��E����NĵNoԢ.�z}M[�0�v�ݤ6�`sp�T�I��o#�yWB�&>rw���V51�2?t#���,�Q�Y'[C�x\Bn��+=֢�H �����~�}CD�ݛB�h�'��Q�1������_��v��Ф�������s37� ,r�^H�r)m����������Ӛ?������>�K���s�nr�޷䣈W�xő��v;���	�h)8�rX��Z��?9��y��U�OX��b��0�F�lF&��	n��X�	W��jt�t�`$#�G߆�	�]����=/�h��ʲ��]��fI[>@Pz?�:!�bF��ڍT\c����
7bm�$2��;��|�/������ș8a�U��U��*)�/���G�B�,uQ�s�H���5T>�5U d��!��Fv��/�0-�"P�{����$� ��6��]B&�u'+��)�����q�X|�Zxo�Ԋj
D��m��L(�`�.V@����5g�_���^�D؟��m���%��g3֛D�H#dWx~h��6ݼf�.\��v�W�c�-��,~�EU�>�WWC��0N0Co�sx��l���f�l}rI\b�0�l�,�&�AW�'�/`՛� {�*o�i 9��8j�����_�a��lJ+U���K&:���VA���<�S�lҴgB��Ƨ���l���K��k���N~y��D��5 W����6I}�@i�y�x�xŠ_ �L��x�^�U��˨?��HB�+zs{��̓�@�����~Y���c.2��Y���UllY��s���զS�<��=��xt�"c3����i��^Ƌ�l.�'�@T�p�������-|gެ1ߵ�"'��)n��V9�k�E�@d~��Z%4�=��_��2[��?"?1���Xy�1#����~j);�nV�6���ߎ&�H� ��r$��X?�����'�qҚ���v1����e��Ԙ�_��N�Ժ²�����[�@��~��~�s����%/���0\4m���C��khb�*x5�pR��	�י;�]wp_4h���(��VZ�-��������3G���-�'�`�*�(/W�:�J7�2�\�������[�<ֽ0w^�E�`j����랬��t��G��������d��p�yy�aS1h�_b|�ox��;t5�PE�n>��Sx{p�j ������V����f�5���ss���'��i��`��py�B��41�	oX;%�A������֥��I3�I��pv����,w;y{���0L��ؕS����'�w��zWCan�z�B����+�n���Ƒ����6K��=�o�u�Ko�=��k}�����1xq�R?+�E�<��6;���M�������}A���EGe����Ȳ����#������w��m� !A���&���0����z������R���b'�ͺr,m�8-s�������b��&��6��m��#��iA՛!>�D��mL�9�3��h"�Z��.E����n�����Ƀ�����e��^m̀h�0C����yB�G������h��q�v��q��ĩa6ԥ"u	�8-�A�rv��x�X�+ewE��W�����^�������<|'k�����%u��λ&i寂T�
{���Z���ƭӉ�23�\���jK����P����"�c�dR/=�ߜ�6T�6����$�%���ɔ���*���Aa��pY�!�!��)�K�ϟo=-bwf|�t��n�᭦�α���<��k�ʱ�c�x,��-��1'�����Ԍٴhu��G|�����ՙ>�>�A���h��FG�[���IsC���7��S�飭�ed�e��=!:?��躛�)����C�w�5u�m�Z�V�R"�
��"#�
����
**� �VA@��T�2e�A�=��V�����|���}��O��Gr�{\�u_�sN�3N_�M�'�[����Gܶ�ͤ��b �M�����Q���Ƀ�C��ov!��g�yt}�Q�sxo�oQ��;�˰���G�������8��uKFS;S[}����(ë�fPh���D��/��e��g^5�5.J3K�~�AP��P3�1��Q���gY2UVkZ�5N�G=8�>��]TXK|<��g}
�B}z$��R��{T)
|��7��\��o��k��-�c�7���P
j���[��vd.����~��֤��?����H1����2���8���]�kc&dwg����O8�?�:�(��/����T���v����7�����?Ӕn�nu�3<z7�SK�O'ӗ�"��&3���l�/�j���ƺO�k�@���'(��\U�
4W#	T���Mx�g�|zj��4uR�im���=�/�O�Ĩ+�}WMb,=n������*f&y=ƒ�]�."��o�ٽ��"�"٣����e�ј>�UU��'��o�k>0[�,8>�Rx�z�z�� �3v9�>:yu��|�.�]0yw��Mn�\�����X�7@}Oؖ��ʢ�?l��ڷ���e~���+4
�|ha>�Ac}�f�"��A����+`�_�:l�H'�'*�?K�GW����ڨq�"T��ff�F�*�.$.���a���?+nL5�p�OɌ��U�"�V!q�_O�����g����?��
v�����a��p���� 7��V�s�
�{������XI<�_�Q��-�)0���*Q��W�{��7�N�H��QP����(\�N.p�2���9����i�WiX@�6n�U��t:�BN�N��}�a��ċ�z��=�6�`��Z����|���&���k��`��ƞ��N�<N	��1�د�~��B9lDN�q�W��%�嬠A�e��qD�~��ÖW����[���F�\
���k���D���5������11�Ig������|�4J=�!*� h�IU�c���Q��4�B�`9���,��*�"�=�C�5,=c~[#���r�Av�r�t��-CPJ�n�!cqjG���o6�dV�D%���'���e���G�9����ŵ�	d>��~�0�u��k�M�Ŧ]]Z1��t@�$�8��Q}/�\'��ɵ�� ���aa�S��#�I�kl`���A�&���E��bY��
x�#�Dgǩ	�98+X�6=l>p�8�`�{�뾕3���m��R���AD�}˙��4)DP<Iy��S�W9n�����J�o0��4u�M�PC��|r��3l��br9�{I�	��·�~�Č����O�����HO�	TC�>y�o 2�X�����(|��W*/��T���/�����k2����J�T�=���m=[Hf�NйVX����a�9���	��"�]Y��o��{��UJ0%6C'�������>>z�S͇?x�fg�z����}�"�g~է�οd�;��>��( ���3��R�PC���~p�t����T�,9�^�}��B�x�Rp���.k-֐����:�m�;� �l?�600PI��d����_c���Ke�c뱜�����z�<@��[�d�`J�1Pʞ�cpG��8!A�+9��J�n-�a��g
��9g�jT<��U�_r Z���e�����+ފ�?�S�ey����X�|T}2g⦱Z���ӗ+�(tk�,�hc"��y��>��G�{Sxs��(�]4yc�;�>C��w�=P���p�93$RX_E�:r���+v����J!��wx_��آF���;X��D�/�����o�%U�4�,�v�����v��eņ7�x�QL�	��~\ �AP&��&gv�e��1��ێ�n*6�ԯ��������a��[��{w�<t�<ZnL}��|=y��Y�	~$��\�����+t"� 3X�;M�m��t;��7jS)y�v�k�S9q{-% �����g�}d�,���[��6��:P>]/�}X�P#f�V�4�ZL+X��w���� .�&�%�C�����W=UIp~�	�+k��N�I"ӆ��/˙ga)_YL���i�������s��u9A�Q�sG�7�s�at�{�&G&&�10������{��,@�����?�~��Fd�b��ẀPT�P3����{���շ�Ru�|��gzh2�,1rY5q"��M�t����Q&~�ʯ&��B���~���g�>�̇O��e}V�2'�YW�A�{���{�`ZI�F��ӂϢ��U����ؑ
�*�Ƣ�n^���~wh*��9��_��}���������o��ć�jnmF��:�D|��We
�D�P��w��:��*"�U��2��%���U�nc�MK�ح��^�q��I���uG� �^�hX+�a�������]E��$��<�6�R�ɫGz���3|���K������֯��`=]��mD���i�b%�ͩJe���rM��Q=ޅ�;Fc	M��kgO������QK��d�J�X/��x�P�D������T,/�*���%H�ϰS1?�wpC���c$��.Z5��F��k��7^0z�@��i��� �m�ZOH�s���<�do'H�8�{h
�+L���l"���UD��mp��w~�dT>O���}��΀�t%���附���Z{���Le����w�t��e��@3?S��U+KtG��jHY-���ihHb�c�Y�#�ذ#,�/i�v��و4�\ .�z�uE�
��q���T��v��i���}�q>���5Ųg�� ��Un쫎]��l$(ץ����:(�2q�.�?�D��	{7U�Yļjji^ș�i���é��s�)M����M�f�O��}`��܀r���~�p���#ܩS�_B�'�B.�:���:h���rz�P�3r}��Y��2��)��vJ��ЇVǹ�ꅺr/�Q��ca�o�ԙ�M4���ҝ���y�wʧ�f��֖�R���S�^�%<�
�"��v���}�T���q#�5���(�Gk��RB�ڪ���k�>�O�� ���f�	u������t����ky|@A�U>�IWe�5�b��JJ,�j]9�$�w�#�6��2J�Ŏ80�#ԋH��"���%�B�P���6���U�J9(d�˱�V����6�}�.7�MJw<�3c�I�9rKպ|FWz��wh�Ц���+�Ğ�i��
�toF��*�W�ڴ�@@�F&��aT-V�h�!(%��X9�lp���I��l��"�f��~3Z�UM��%4�(���:��N>=�h��{QA�Z�K�8���0�x�A[��d�(��K�>�Ğ�)�˛�t]�,԰��@�˝��~ܒ0�p��%gil�]C�Q1p�Ɇ�F�k��H"�g�%�!"��N���+�U����D߉U�^�yAk�}΁�z�dj���F~�O���\���!^u�'��0���^Ԓ�r�� g�8�9^UEq�D�r������
����K���<A��CWA4��ze 0Y��zw�fZ�
����[��c}�&�[JR�Ry#s���s��w����4��4�S��H�t�U����	87ŗ����c�'<�Yj?���o�;Eo�O@�P��z�Y����,q� nY�ǘ��ۯ�l���kM�(P߰�����d� ���u�K�]d��Ʉg`���I�2��u�m��O���r�py�t�#��ˇT�=T���~���Ь��?'�bϧ]��:�� W�)V���f�5�����cxfbe���)��Q���˩�Y�8&�a|��o\��2f4
|�,�	uǘg%f+M�[Z9#i �Qvy2��䦕b��:A�`?����ѝLW��(�K����`�>�����uos�,}�܊zHM�� rE��ruHN�2ٔ�n�y<��l"_��xd�S�����W��=�͎�@YC�ƨ>�wl(��<��Z����Z,���qA�����Pp[E�h9�[Y  �O�����fq���{$�����r��|G�U�R��z���p���a̕A�+u<yF�|�e�imoF��9�0W��]9v�'=�Szp�~�JG��e�X[���;��HFi0��C 5��.�$�	����a�<�?�~ �J�W�8t���SU�������H�W�<kӌH>V�� F��U�X'����qb��]��w#�z@��f5�����%���{��O��d�ꛆyL��ZD�u|����,'I��0�l�q,F�2Û�u ��&���kyR�ֲ�ˡ�2@j6s�r`��ﻻ�z���,a�4u�<�E��E����]��:R2:M���]]JN\��I�h���^�'�a}����ac*z���oMmq.�H73�j����dv�)l����?,p��k�o%;,͊��Sb����p�U�G��r��&~�Jl����G?�D���W0hvs��p�&�E#��rh.�%�g;�`�'^=�;�U1�����Ϩ�-Pz�7=� >�d��A��c|ZB��I�e`����uD�/�����JƼȜ�VO�U[`���	7B��Oϸ�^Y�*I��}w�޿����޴����&��>*�ޖ��;oI��+�UW{-L��`��D~~+�R�~D_է�	�'��E7���[�*�j�˧5=��R�q8��Sl�zOĄ�wk����5"c���y��-�#o���C>�|��|[�����[F��䅓��I��r�jߏ4�Ӿr=KB�8P���S�I�h"�4�����V�MU��c�;��3�/q�9��_ }|#�%���䷩�8���^���G�b$ac���rN��RZ��L`M����dUTx���֐��R���JQ�D&c/gtٷn/N<g�D�e�҈��{�Ti�wM�! ��GU��9V�ڪDU>#%#
��9�$�暛�D�XZ�����^P}PCWHw�n��Q��|����l�Vp�)���P���{d�!�'��y<R7Υ�E"m��]-����t�o>�]gt3_ڛX,�@
��������[�ڨ��(��(à6a ٝ߯���]e5[�"w�#&���OX�5Erͽ�C N�Y�g���]H�������Kɟ��+W� o{�hY��Qb]�a���/c�~����,s<4�1!�9){8	��YoE>r�n���T�����zeJB�p��#&ng뢈�v�q��]�����z�-��Sg��iBl�"�Q@)���gU��f$���}w_��Ŧ��(b��g�H�X�%���V���@�7��Jq�N������%A����u�2�F��+�+|`?���~ĿN�4��5 hb���(���^���h�Eߡ�\3�LS�3�|�?o�!z���h�H��.?���7AuwX�#NV�Y�,���|�0��	˪��Ikau��������#A��O�d�y�+,]S^]a�%y�&�)R2�z�r�(�#����Z� ���kA#��m��BC%�2�V��P/�X�t�l��O�G��sE�Xye���ҁ��Ȏ���$�i��Ώr=i�{'��v�Q#
7Y��:w�cѧ���8�=b��\^�-(um�std7uA1��d��t�MVD_�N+�Nq���k���XϖL�q�S�8�>�,:�cߥI��N��Q�
������+C}gT�|i1���|5@��D����:��#�w﹙z�!�*�*��`�H��x[��o]�|���l�
�+�!n�� �{B�|I��Q��@$S[h�fh[�ai�>���B���:���u[a�)���rh��L�6ϭ��9���i�u�7�+�G6j��B�
�+`���-2��W�����z���؁B���lp%R���>,L>�U��琹�윌��(hu�4��툶�ӕ>2bҁɯ��.�68f���>����gͯ�[۶�A	�]�ĐGk����\�p#u��Q�D? y�_g��ܖ?�����(@R�i�k�l
5��
�
c+����|Ŀw�P}jv#�U�7���m���/w7�q&W���M q g�Ip� �OcC��go��V���	cum-��$��K������8{.�F�����L�hϺmk�8X����چ�+Jq��|�O��D a��6Y=ۆd�?���	�.����
�����}��u�C�3�N�	����C�
y9p��þŎ$ܯ2��=��J�fK�di^����ƹ�c��� 	X��W�o,�X��ڝBF�N��K�x�|�X�<&��>!�_��+�b?�.~WZ��N\���6�ͬZ���`$�ѹ�X��4�(�X;�����B�`&��N;��^�acԡ.�Z&��������Z��T��dO��2�Iu��<��h�S۲ᡸC�-���g8q�M8��w���΃�0���+%�c�����e �V��vm�[9�����i������Q�����V�I��� �w�9�s���˃D�����������]�c����?���e�����c����dtO��:o#��	�z�������JQ8�'IGe꿙$v*.a�x����Z����D��:L�-+ϸ��ʹ�l�LPp)w�	{)ly'�/��C��"e���797�/�N�W(߰:��u@P��h^��@��]g�7�Đ�9ŭyQ|�f���sKM4M��w��t�n는��݌Y�-o��F�r��p��N�f���^����������7�8�J�IkcۂD��������"��}���-R���FCC(�$0���\�_6�*~'zs��n �/q��̣���?T~��E�UD�"�>Jt�?����L�4�nuT?~ ��Ð^���u_�Y�,��2:�uѦ6�+4 L�,�h��y���IM�Ҫ�w����]%���c�8�,�ןl�O~1r��e��L�方��{t���w�Ƿ��d7����X����8u�m[/Aҧ����1*g}���X��M��䳖�uq��H�}7j�/����Y͗�UE/h8|�0��&��l���eh%�����DϾ('3���������Y�u��1ߞ�h,e�����G�HN���#�gá�h'��� ]������h�Z8�Z2�飄�	����[�<jd�>���>����t
>�v_��U��:7�G��Q�o���c�����]N�R_�˼�r�:�Rfc�qaywM�կ��T��Jz�˖I���(�l��� ���%8�n]h�lli��5����A��;�?+�������O��m���VϬ<�N>�ݼn�{��-m��̞��o+��R����VA���WxP���f��cS
qu����8��U�,��^�4�f�x� �-N���������\��[�@��L��i�M���V�B\�no�"c}!k���5^H�ɪ� �F��-8K���>J�W����y��M�����Erݷ	H�|���Co�}�rK[�����(*��#�dAh���s-+�&�F4�X�y��NB5Px
�Dq�'"��?�Gb��L�#����8����΂�J��q�E��� Avj議7xȁ�i�C���a��l���n���g<������#�� �7�%*�0ͽ�[CnKo�+Ă�8�&i��>��M�)�,��m{�-�,��2�$�	&g.�i�0������2&�o6ik(�L���E��d�u����ε�ӑ
��[�<x����s��k��G��cK-X�W��[m�=�2����9P\-�V�� ��Zk��Ҷ�ǯQ��zﰱ���s�q}̡�A�l�JɻV:��0^��X�ndO��6�c�n�1|���e�t$*8��r3!��߲���E{F�l�k#��P{z�:~cN�晙��y4SQ�[I�1�Y�R�m7mo��u�u�RvI�n�U������G7XO��S�B {6�4�L@���nM��m�|���4%Ӗ��h&�4��m��3�.���de���VV{��	�(8���xV.p�")�(�h��e<wX�i���~Y�#8��N�y=86�E����n|�a����������L9��f�I�O_9�
dr��#u��Ļh�����e]r�Gh���2H�G�F���+��!�T��%c�q��ضy�R>�|tۤڗ�v� qX}�4����t����έq��m72S�0WVz�&S��E���2Qܒm�TZ�%l��I���˔�۹}��&e�����d�̒���B��*3�]@��=M!�mK��Ih��qsq#��^�6�h��� R���Q?��i._i��f�}Et@����A ����78C��;�V�b�'��a����`]�*l�9�6�^���k~vP��X��Y�r!N3|��4hMc�̰"M}E�Aػ;b�.���<܉$���x���7�7J�s��n�r�����U8�Z�捣5P��2�V�p�k��N|��N}�J����L��Z�X���6�B������C}���䙊��k�\m~�%O�ȅrO�DʉԆ�;nq������ۍ}�e�m���xb�Ci��`6^��rJ��9y�������,�4��*��ݦ+�հ>���h����/�r�7'a���[	�@�_� {����V1�ݦ�H��/�6���4��o����Fz��j�K[��&���]�#oa�u�����_L�)ڋ�ℨ�������և
n���8���>���!��;�!�嗪Dwo��A����ӷ��b�n����FC2"��t�9���a�0�׼58gZ眈~~�Eҙ3��Zä�I������qI�:,x��>����f�J��>�<7ѓ�Z| 0`$k0؄�˥ �'W���"��+���\S˅g�Fr�-5$��%��#������6f��A���?{�[��e;�Q��0��Z1+�Q�ޭ5x��[�(.z�I'�I#*���*$%ɉ�v�\[}��l��y,$��8�?4v�O&ƽ�p�d�Q�P\�m!#&�T#���	y5�T��.S�Q�0��� 6�E��V�2�?����d~�~��Ȱ��jz����ǯ�XG;z�=z����/�|����qr�S�KTe�8y�����r��l�|�	��:�������M&UU�֐_��3u�U�yY���x�I}ai���h��r���9C٫g(D�m���^��(�u g��y�G#�`�a�S���1^��ȣ�o����8�/��B����2��}^��ϰ��eq�<�����w{���ԴG���=#27�:�57i�v�[/��U��r���з3�׶��Z^��8�[i�U˝��_O�Z��EZ�̭�1Z�Ü:����ۼ����Z
�{��&Q݇����:0f`��X�g�6=W|kr��Dq�Q�^H��\��_��Q��m[U�'���	�O,�Or7�c�����,���/�(:9��ӗ����e�X9�.Y������V
�ܠ�{�wN?\m�Z�w�yp��='9��\��Δ"�_�H^���J�o���fn�61�|].�R���'���n���*KH�¼��jjk�=8��=����S!�k��-[
o35�����}�͠D��ʉ2:ͳ��N�S�N�1����U!x�ݪB��Ҧtc��`��ŧo��A��R^7eۜF>)�u����cKo�zQ�2��P��P� ^N������}�_v���c�[�,�����y�W֚�|iWr�ջ��3޽"'3��KQnS+V����z��J���\�AF��L�٭�l�@.l����ܶ�H/�z�k�loT�X}(D(��#o���Z�~!.��]}���zG�M���|k(������{�����Q��6fd+��3�$Q�����݃$�d��dKЂ"�A��C���c��BE=#[\)12�e.�g����֝;u7Ζo4�`Q�W@)�}���,��u�'q�#��a��[M�3�zȡ(+�6���%�V��Vx;��x��dϠ���o��P���a�.l���?��ۗ.ig	�}g�8kx~&���t�%��֫��lg?�:���jK �^߾�5���r�������b�
�Q@7�N�R��=�
Q,���;��������<�l��ߊ���W��P�,��C����ɓ���&��i�C5^�m��l;�j�C;	fj���@o�'|����2��Zmn��C�H �W���o�$O�sF|��������-1֨�o_�X<f4S�ߡb��ײ�!A���9��S��rԘ��zD$��]��i,��z�4���f����C��Ed/�k�>�-�B2�P�}�Fr��Rm9�x�J��1yW���o�C�J��MѣqK��u�cjPs9'��!\,��_]L�kÃ5��iǾ�@A��&�^kI#r�r���9I��S� �]
���P�j�Y���rtG�.����h�y��Iy����㓇IB�Z;T���S?���BQ�h��h6� ����5qn}�6O����"�;��T٣΀�ɸ/����@���^К�4��yﺏ��ٓ����mL��<����9%�
;;,v����G�!}۽-�L颅��W�/ |�Q�N-�Y���dה��t#��KX�'V.)�c�{�Wdz���%KyJ[���Akcj�J������i������)2�H6��]>��m��${���(��H+̠���Fc�r/s�xIX��L�����ְ�b��D��^�JAf��&�
��������*�O	ޚۿ�+h�4G�Z������i:�6u7��/���M70R2����(p�����B^(�S�q�k��`���Xu q�h��M�/KZ��Q�WG��2��&s�'+�k�ڄ�w�2o���@�/C�����m#�֌��&F�Xi��[���`��fa�um���܅���08:��.?�Z��6L��W@!�j�@����Nd���#�iHh������]��'��@��M�������D1C'k;,�m7����'@<>	&�d}�=^(�U´��"���p�
��:��	�tW[x�z3Y���ff ��PZ⡤��D�B�w��� I��"�j�0�����dݹ:{��:j���������I��_�Mӛy�R|��3t`��X�91<⇳' ����g]00<�Nl�d'��mp���r��?��%乙<�Tzf�๭�V�J9�={>������ ��y'O�j9W�[Şw�������\%A/>u��?�vǻqE�v�Pd��HBWu����YB1t&���]�f/OWcy�ipO�|+��ig��\��"c(-�h/8D�#qʖk1��R���P�HI���u�%�%��!��
��{���)����4��z
<W���f�ڻ��օ�*ۉ��W���7�ꚬ�
��<��'u��k"6w��5��nqg3x������$��*�~�%ry�v2יWq`���څ#�8��7%�U���N�J��3�Y��uy�7kA�#\�R���'꺏���u'+�ߨU6�p�^s�V�E9�L�?�L�"��:x(z���g_�N�<ߛ���'ɿg^�� ��;�'s�n$�W�˽Q��@�$��t�'/�C#��+�k h�=��FsS�k�sAjjf����r]�Кᇠ@�˓Vw�f���z؝i}`��p���ډ8L�NQ-i���,7 \�D�[2Y;tA!�/�4>SV��=h�}®�e��׀�O�-��������w�p ������V��O�[j�L�˄�+����od��F����*�
"o1w��b0�tㅶ���w�/�'�qY~S1q;�u��\ʬ���9��}��+
W���U�/����J�L2�^]�?P����V�Q;��-z��ܲ{�ѹ:���2X�i�
t6���1B�����K���9�}b����%Wj6xw|��m������,�|9Kg�Q�I���4�Q�]�y{ΐ39{�CM�����2�fCґ�d�;dgP�|�B�H�!-<������g���45i�l��H�nri������׀g1U0i��&��N�;��6�&C)�]�ֵ'K��n�Љ�)�S��T�c"&>��|�@�qe�,Aj�kC��/_fk���6oT�9����M�A����RT�_�?xvLxӸ_���hs��ݻE�������T+�Z'߾v�|����Wu�2N�ޓ�5+�a��zծ�lb��G|L �;�xEvǳ�n�`�0l�ibD�o�{)w�`��c~���kd���t����5�y���D��)�g�����[�|�j��`_��D��MK{���eV�H#Y�s��.�}`���.�b%F-����h��� ��Y��('�p	��T�i��� ���@%�>��~٦�����y܊�r�r�N]t���0Hcqv���߈ͦ�E�^,��SR�xW�Q��o�xn��9�c�tA��lQ
�2)��=B�1��B�|Z��f��\~{D�we_��b���XK�ڴD��ֿW>]���>1y��_��2Z�˚����4˷�'������QC�������I��"��ٻ�}�	�>jy�ڟv��ǽz�7��<@]\�O�KW?
��%+<QN�V柚�1:)l��7����ӶO�Y8��,ᩎA���	5'm��ƾ�ׯ�t>������ӭ��Ԋ)�2�����z�Pk>�^�ͨҞ��\Z���ȔOQ��۾kw��$" 0�)�|f$^*�7t.����z�A�Hd�����m4�X߯x�TL���!��I��|�^2��p�����%��vu)x$�|ɦz^���{�\��N��@�u�t�o�������*�"��'U��9t ��5�븷�)�@�@Al��	�mओ���}���*U�5����N�g�Cwl��ulZ
I�c�Dc�(;%�N������i����"��JX����L�@�<�@Z;us�[���E6C �2kq����$+�(�ߠӓ�gH�1���"Xk�MuN�p�&�y��äD?��.'�93�x��)�Z�WnL�M�=wO{}dtz ��d!�y��Fy�r�w�̬��9����E�V���`&&k�p$�c��=�eN�0c�\��s�v��"����/#.~l�ư�� m��B?�3�4k��ٵW���@�x;��8u��ۆA�9XA�W�n��C+�t���>��z��bw3Q��w�a��fQ����zd4|%�7�Cg-�iB_�n��Y�cd b�2�=7k��y����b���AjՈ����T��5�Ơ<��|C�!gNV��5qWï8�s������A�!R�cz3)�o�C�B�KX0owN�(��×��T��{�AK�Åsg����������VI��)#&�V��Z6�[�u�KB!N�i`E1Ndj�$��p��<8w7���Ѳ�^�c~�b�=�WB_]�'���KJ:��.h��ɘi�<���^0<k2��$	Q8u8�϶J��*��|�B����ň�fö��*�����	�/_>��ج*�兔�xa����������7)*�o4p-�|xȱm�����d����H"����@c�u���1��~�x�haXDd�(tZS�>X�?�Zƞ5V|�.:��Gւ�@N��`��p���E��8�ۓ��$�=�ȁ7�q���V��R��(�BK-���C��o~�6Ԝ5$빼����\�0�	9xt�}}�u�u��A%���L���	,�<*�_1�ѽ��hCW�>�<�@���B�T�=��S�-�9J|�MW���ct�OZ��m��������ʒ��>�l�k3/��t���M.�FJ��#�4��
=Q����-����:�Al���W�h�@,�l��aZ�����ƃIX��Sj"i\�NS��%O�rDߛ1�5	뼳 �ZC9�4<4z���r}�ū悎�B>��� �$�a�>E�˴�ٝ&�IPeiyR3au�C6���w�=m?'�8	0��|����͌�R(��RSjQ����vJ"ynz�Z��ۜ���CC~���-��%��C���-ȸ(�P��l�ffGDP��UMɔ���4
A�d�
W�4s���Ӎ���@�*.G�h� 4�T/@\�jX��vnz����C��U�S#��>þ��Q;�j��> �V�mW�aF������7��uG���3���B~�b{�Oh3ӣ?��r�DUD8=
j�倴)+�$Z��w��c�zC�8�aF�'��R���r=wNO:B���E����G�z� G|j��i�{Zˬv�rQ�N���nH	���w36��Os	���Qj6E���	*��i�sj�F�F��{Mߤt?V�#-����Vu~LEX!�]-����w/Fʾ�$�t�bR%��l����)�w0���	�[�e�F`S��C�Jtα,K�S��B6���fJ�����_�TF[_%XX�!���>:z�GlE"P-�	��c�ݥ�v������?�� ˢ�R{���MM�]2Q^�G5t�i !�j�f�d�1 ��5-�6��������֪��zX�Ȍt��#���v2�G�x��R�8�b>`����Tp�C��gdqs#���%�M�����ʆ�c[��F�MoK!�[(��
T���H�����o�&6�1�*}�8��b�pV�q��Mk�V X�_���U��:��F@�~~�cԛ�����8�m!B��x�N�%��I�ii�Ii�h����1��eF�~(�h����hϤ�W;5Ly�E�􈩻4$�9��M��hK=E�NSuAH����-]�α�~'�qx�U�A����t�{�!�)��R�6�x���V�ӌ��-NSZ�Q����ٟ5btN�o�pČi6�gb D{�����<��Ԗ����I�53�9�`��lAk� ���7���@�(GI�3����O@��C`Z<T�r2�,>��$�<`a��d�h����K�]1�*�C\�����*ņW{S\� LGv�Ak��.�2`Ā��~pO�$�,O�ʄ�A�GdXyعk�Pn�܀�#]�9���٢'5�'��6��	|B;$J�t�b˺��,T���#,ĞL�.�*w�P?j��DQ8�v�O���3ɋ��t�
5������x)i���~&�&G�N�0M�z�z=���Q ��:�"TC�9P)��������c�C�T�z��~�����T=\
��Wݲn�:J6��q'�mZh ���{Z��Gߡ���ꈯP��#�S��4�ۥV%�@ o��yO�qxZU`j0���h['eX��+=v-��zo���b�P5�͈��Ix�ă�R��'Fr��\��V>�	���ǎ��5�|ݒִ�"q8�43�0�G^g�$q�zq�|��}G��>����Ӎh�����4�J��P˂��K �>��n!.Ƒ����i�L̟��#�3䃮ټY��C"�D`��!NQ�)������Ѣ$5�HQr��ߟ�(}O��NZ`��]��|t����1Ϩ(��n�~�jA�0ҫ�2� �U��� }y�G�&�;�#6�8	(�[�ux�+)�T�>�$�+7U�d/P�N���>���a���V`DE����ݼ ���Bph���z~����3��U�1,�w��S���~�<S�~�O�#5�m���N
dm�����	4�獀n$�5u4�tt�Rz�5�S5�k|��&��ϖ$1R�O%e�<��D�G�vᗦ_<2_5w�#�g ��ϴR��̻�,R'��,�Z��d��J��H�����pqf$�7�(�&�X�^D�m:zCX�γ3�(Q��(�l�/i3�~��ZS1-E�V8P���r���$��BտOwo:l�D�`�R�ʡ|�Ł�T�1���ׅh9��E��e���]5�ħ#�r�O��{S�v)|�RWs��_����	/��Л~k�����u@���:�UCۈn[�Ղ��F��ʪ.4JGX̩ԥ�d�+��9�h�3�R�hA�vSN�eΎ`l�ڭC��N�tCO5��Ε"�=@ԤE���7?��H ���k���!p�x��Z	�%�7/�6e[
gīU}u���?�Y5���R�Ju����c|�*-�?�g�+�'��R����Y�ow/�-�~�Ԑ�7�X9��q˥E��XaU��0�J{n�3���t?��'oI�ݖf=���Ԫv�%(*��Wx^��z���ϓ�tnI����įCP�ҡUU����2��)Yaxd�_A��e�\��Q�	/>`���М}aKMհv�!i�e`��#(a�' ���+�U�I�)�a_L氚��Y/܍���?�z�`����x�0v��ǰim���ds�\[ �SL#*}ӱ9m'��x��ؤ���@u�OZ�n�����s�_ֺZ�땽=9���Bn�������+�FA�궝�٭�{��6ջ4�I�8�Rd�u
 �Aٽ�� �AF�5�Yt�>���z�R?b�y�\D��z�  ���ڧ?��H�K�H�٩�}~K�4�|B�O�}� u	�_yC�M��"(Nc��о����:FZ�����߹�A�Z�E��[�%J������C�Z1��!�� ʸ�Ȕ��'�#����.L�%���{a��nAǳZ�٧����4c�@�%�.6&+�} �Z����h���"����_H��%�x���2bRE�&Tӭ��#�3lL�pq�D)[���n|�m�ן*���XR �}���=��s��R:p�^^����̽���p�{A�F��n�'৬2`�����B��i�҃��y�׽ �����Rb�D	�Rŝ��SuKǕMf��"���I|=��%X�]�L���İ�т<�ه��c��(6�"��.�ߡN���\�cX�MJ��B��55B�d\�y�a��WZ(��{�z� �a1���9��U?t8��=G�xk��ZG�:�X�.T���r��KkR>C�4)]ТA�P�u�4�9i��i�����Ǫ�5�15�`5�g8P��
v0�8T�]@�#�����3i�3�/K���:��PLEE���ao�=;��/> U?$ט�d���j�v����H���K��gl�]�h�ŶwYaVq��bү���Q��/�Ɯ,뒘F�D�Q�_
V�%���W"dwcJ�Ӌ��$\�߽"8uK��bPū�1W"375V�"�VA$L-�1(�[ɢ���r^舻j�4�ܗ����͍9�7����\Tt�\��FU��W��̝�s.�3�w1 �z���J5�W��L��W߶$Y'���{�C���)�^x��W������A?~����)� 'Ѕ�)��Bω�K�j�qp����tD�0NiÑ~��^�O���w�G���m�Ì�R�~�D��S����ғ�ɛ��f��oA��n�&��9ո�k�Q�<��o��¬��{i��q�*��H3�EI�$!J)[�����Y�K�	�s�2�`{/����
#}J3�83rM_Z's���HJD;k��HH���HQ���t�!A���ם��C�g(�F��>���S��Ӽ-iZ�pm���� ����@(��MU�����]�����)��^�e�"��]l+:�u���.�{Z�P$���Tl������aM]��hZ[m��� 2���Њb+�2*�(c�A�[��(SdT1PQ�BPQ�QE�0	B ��a��O����������}�+�Yg�5|�g���I��?�m���4F>%��ܜH��=�Bh;�ejmY}����7/��O�[q�됪��
n�lP�ԉS��m�h��ڛ]�7w�dk��׽|\貴�Yd��U�@���-j��C�e⠅�й_u�|28�|y��S�}s2���smk���e��:�rvHTy��g=�/��(�ʬ��OŊ.�kyw�ls<ӫ��/m͇c�Hq�j�EG�Z���lֽ2'��o� (;:b�� k�p��@�vߏ9�#G��rx�6��	=l�B�'��'aS����h������8�s���M��`hQ��J6�J�J)�1��l�D��9�c�qv�L�����������ϭ�/v�/�r>��i����9�F���bi��%�zƙi	�������f�����,fgm��F{4�[�$����wD��ԭ-j�Vv|��\��ݦ��.WC[���y\��[��_p�*߼��ě-S�����ܤJդ-�E[��Dq�X>����L�;�ې��W�<N� ��U�yZeg�ޕC�[�
����T̏���7��h�f?3-|��@�~뒔v���L����e�s��=��1�{J�Y��U��AZ�OK`��0�i��EO^�������l_�4���ͻ��E
:m����s'ֆ������ZG�$fc����O}��{y1)\�%��{0|��&�`�y��Wɜ��6�:�z���d�o�8s��0k�k2��x��s�ܵ����6-Ky� ;4SS&���,�^殝/L�����{�%jߩ-�a�u:��ȑm�ʛ♃>���9���������^%����T.���,¿O0�;���Ж��33EPĞ柯z<?�2�=s���v�Ѱ��<U��"��Q*tXlp�+۫��4?�!D�[�6�Ŗ**�}_w��۝��RO�ދ�i~I?d�Ie��~v[2כ:��O��i{-�Ś���}i����u��p �_כk�����O=����/�&hs�ν���}jA��p��@Q�v~j��h�1d(9�;�nBU[��T���nm9��7��`���#�ˬ��]��׾�������pq�Hv�ýYy�����	�l�W.�E�8;cWMҽ�of�w	9{~�DŰDf��~r�~��!��y�����u	�Ԥo�b�;͹{�_�7r��{ʾ.����V��Z�t���]��u]4�^q�`70λ�og]_tF������Ӆ<��;�.�m[5�8޽'ӣ��2���o�.O�jf�0P��)Ӎ���C��'�L�~j(k�}�}�77�:ER���~���;�s�����ǜTr䷩��F\J�T�ޮ�����-yS3@���+cͮ��S�N�8�q	���5{�G�Ή�,J���4�j�T�v�"��U���xV ��N
\���R��&l(��Lz�hUJ��#���;��O�+�3U��Q��K�yX�|���!-�
�ڱ�'jS�g9���>�{��̥v��q�J����Ɨ8�֮��`���_u��d��>���gpx��+���\�l٫޷��dC��EL��5������g�n�����/��uM��ph,�S���+o�B����qM���������vA�o�dR��K��)���;�|���t?Ns)���p���;.<��z/��i.{�+�}y;�7���~����<�bx�^�H���r]����.e!����Z��4�8�^�tk�I��r��v����mZ��z�K�ք�}ג<���潡Nm/G��-ͷ��o	���r��hΖr�K>o�s��%�ʉ��-�Z�g��l��q�~�K��ŭ6���s���Gj؄����)I���Ι����)9�)<14��z���ӷ��}i����]y����H�H`^H_E��D[H_�&
�1���Ɉ��iZ�;��o��~%v#ʚ�$� Mя�2����oP��m���K��\���/�~��˥�w/��qBO,P��d��OU��|;���Ҕ/��������Wj�7�Y��/���՗W_^}y��՗W_^}y��՗W_^}y��՗W��yu�w.dK!GdJMA�KS��{�2O���m��K���.�k�����?=PY~�ǻ������!L�����wk�����k����oB~:�����L���Y�~A�����I�Vao˴�̷Y)�)m`�]��qj����}y�˛_����7�����/o�?��?���&?�3��x�3��?z1��]�$��#����X�/o�������k>3OE)�-z"���g�������շc���|֧zr�����8E|�Siy�E�vI ��	������2�DԾI\JO�<���k9t�,y�����p�h���s���Ѓ?�Q�"��C�R"�PI�\6�(�<"�=���g��ѣס��m����z��OD��&+?�<5'���[Lb���;i��Į[HE7�3{S�<:�^���i��m޼9+��f�\��Ku�&Bۜ����N�/�8�$C<xO	]�?���"7��\��g%2�Se��hk2�������n"��ۻnjj�[�siR�C޶�:2N�Nh�:�?��c����+n�W��}p�$�������������Θ�����T/
]7O����p�4鈕���F&��@�/��Z�-K7K�}��.iߖ��Hj �t�M��;c�*X�l�~�\S���ay\$���br���w�����c�}"�1A���8�����pKb�[�1�R��M���J�}��t����oi$jW���g�E˒���^��[D��Ik�=������AcHl��U�Ħ![E�hS���h���2�g��y�s�Qe]�(hI�1�1�q?7���W�g�Æ�>��W�|��pV���^!�m���yMϠ��իW���5�˰�+z����n&,>D���FE2�M�pd	s��1s>���<���tK�pw�@ø����4C^[�*�~ല� ��Pu��}������"�-5 D+w�6T���X9�����ACiP���;88l9ED7�w9,[�E��E��2\�Y�-�sr�ख़,~�DTم[��[0V=K���z?`�}u������-*��*�ΰ�.Y�c�+�M���R����g���g��/��u�~P�囦�2D�	=��,�4%x#��f�<�W�5�K�|�2�y�񨻅��s��!�_�f���A�`�/iPAN�^��ж���$B~��P�/o��L �B�b�m�&��q[kk�E�. �,y%z��U<Wy}�3d��eFKK�VQQ��	�����p���_^0��C:�W�V��߫��<�E �Й�}3)��?/ ���\ ��2m�֣p��D�U��aq%Ae���8����!e���A)nO��2÷~z�����������/�C�e�9ro���x;��t�ޞ�@�{���M�Y,��k��̹�*/J%l����D�����nT�Bui�Hӂ��|Ցp;&���KH% ����ew�SN�*����-(��!��K��Nu���.#c
p�uIII�	i���pDn;�&�Zl�i�71�NH�W�~���l HЍՓil�v))/��B�4���(�[JDK[\���m�oVf���3_��	8 �ն����7�.�$PR�����ϻu+���D�)�%�
�]�?6��;*�T�\��>��!@�CDn)-����@0����gW�^m*��,�#h)����p��❽3sD����Ÿ61+�|�/%�8�ŏ�E�QT�B�܎)� H�{co�-�%�����'r��3X�O���(77^� +��řC���g?��&�q��DW��g@��h�P9�)�-3v{�;�mZ��v{5튗�ci���UQe�D�7^ěj��ڝ���`V���Mgl�WDk��R�j�cuzL1,�+KO��j��}R��g��sZ���ۏ�22�#
5�!�w)� en(R��f��Гu�?��x{-~�?m,�v�l���b���p����ɪ�ʁ_��|�r|%���&�}b;����:X�ܮ��y'h�_�݉���yB�(�����񴰘G&6�+���,�!B`c$r��Q�W��Zʒ�y �bD���V��+?��͡������7),) Ȋ�*{	h?4��$���o�=+���޶!�o��8j��k�!��W���S�� �} ��[��m�����
kjfP����x�X�;��Yb;����I/@$���.^�i�A)��scN����̘9������"D�_���9���/�-�R�[��r]l +#rǵ�^5)�!�V�,_y	�L�������N��>��ծ����;�-h=�}�X�R��x�Xg@4Ʉ�N���X��!��*��M���DsCh�^�Kܜy�Z	r�$�4J����B�22vh�g����U�"Q;��X%��5��AU�e�9)�D�� ��k >�����z�F�N��u0��B;���� �ʄӕqT  ˣ�v�yg���"�Qɋ�:��ٔ�Q�E��c�hY3;�n~�F�^�<9��K��4��u��E+�5�5�u�����)p�d�M�)��׳�3��Aa��W���5���H=7������4�؝�O��>}*SUQI�D��a��iYY��tT⨶��g�H���jK"����f�0��P�ξl�΍k���y@d�|�ȉ�_���IM��=k�H�r,��	<:�<�,9{$"}S�����+-a�6���Y`�^���X���
k^0�x��#��0�1�����C
I�~,�l�%�
���n��	E��Ak��1Z� g�.�����PbČD�4%����G��NĮ}{�X�����y��%�E|N�l%�"�)���Tu��ح�|�O��bQ���Ot������������c�&��?$���[��XX�D �WOں������?� ���YS��3*+�EK��� *+1**�sx�$���&Q+��2�$�W���i�풱���ʽ�!���^�F)�����m�P��u��G�$�"#��+��(���BX�$��>�z�{� K�� ����	�BV�j��ت� x�2��#@Q�o����`e����xG�:�Y�Jeü��	է�#x[K�6�.�>S��X��m��$���E��%$�猱�����ߟY�C8���ХK9|F�j�@~˽�$,
;������l�M|W׿�.�������&�A}����زjϞ��2���p�a}i=	c��o�v��>�X�ϙ7I��Ą�QE�٩��k1���oD�w$�͵Khx�Oi?��ϟ�8yYY��;�x�}#3p}�J�tn}X�k�����п��HƺW�Q�_��%���)�������f:���)I���������r���LE�!Z){��p�X�_�r`)��4T4�������������K�u�@9�U�dm�(�`��i��4RY ��3ǛR~�ʙ�����ދ�p���x�;�)3��,�KU���@`#
��ƅ"��}a��^��˭_Q��3g΍�V����~UT�&̰�> �q&����7n���,o�Q�o�3p(ח��Z�c,�E�^��x�ňr b��m��>h��]	����0k �V����y.�?6���޵�n��૓����y������0�	r�.,�Z^^�.��������l�v��/�����	��e�a��v���(h�\%o��9ɧz�����(���tJYRkZ�1H��j������9 $JPe?pL�M�@�_@�\� ��6[;9���k
�D�Q���3snu�����%b#i��c|�q�G� f�N���sXfN[�~���B�� �JtV���|N��q�?9�xɥ�˨�p�v���'�@ǟ"��V����ʃ�1��· $H���k�5�U�s�>�l��Ǌ�8B�K�^z!%�!vV���BA�#h�^�i:���s��5Jr��_�e�X��!E�w�Ct��t���:��1]x'����8w�1>�:r
m�*��x��/�BK���KIl0M~��f���	+�x��g	��o�S����	cbtS�'_+�!��$^i#3fsH�;���j��b5J��Ή���"�C(|��fl��׏�:�DԠ�?>M����Ud�U�!>G�'3�x2,�� 2��!S������W��Y�X�V��X*�9!�)[p��ݡ�i�SB�YgB��8����WCͯ|��ٳ�V;��2�xGGo���ԑi���d��J?R�� ����2s�B/Y��s����y�JW�X�?x1'M�T!$�m� ߬A��O���y��R�f���ި!���z���Q�C*�i�A������'�S-}m}�"��B��=���<U��o�
���ȡ ��Y�F���h�x�3/4�g'�Xi)(SF+�F�K�ĩ��8����  �`���Ϗ=��%�{}�@~;-X��������
iT���2��]��cn.䭓��ݲ�-PMޢ Ʃb��Os�i��
C��|���\& (���6�*r�m�Q讁�:-���9id��"����w� ���X�7ۇ��كB�1%�J"�g��R��:	�yj�T�Yy �]��
��$��	5�9���J�1Cyk��;�y�o"�M��Ӵ�p�]d��9���O�рG�'I8�I�-��A�J�`2���ƣ���۱�L+�?��t������)۴�u?GE�q@r�¡0F�K��y0�"<ŭ �13�ʼ��k�Sf���p���b�#+q��r�� TZ�f�O��v� ���3sn��\�Y� �.����s���[PxӮc�\j���RԐxPN��Z�k 2uE�\��v�VE�vKu(6�z:��F'���L}�WD���l�Ӝ;Ϙ8�,��{���
�����o���ݪ Oh�u�^�n��O�'x��}NA�~ϤAM��7��� 8Ib8-{Թ�b��c�SE2"9	-�=p��
_
�/��4���-���E~�\�Y&xdV����"
Et9��^��Y�e�u*��6�Z�	������j�vN�0J���g=<F���kP��b;�LM2&F�C/�����	��6�D��{D$T�
:��#�i�s��Ȣ a[�wk-��?c[�#�5�+�!q0��������$����o��.2&����?\�z�汧��~�ƣ	��b�K�H!@%��$3�>&�X��fnȼ���IǍ���ޭ+�k'���S�ⱄЩv���HF!(J}�GǾV�ZM��>x�ђ��;��~�Qil��1,|�����`$�u�K򮙹�'��J�?∝�{$I킶m���`����#wza��~�}�&	�����W�q�S8�j�8�V��S=�y�vd�|�d�$2��̢�R]�cP(u��|����'�q�c��g\uYcӳ!��)����Og�+n�ZT�_v6�%M��Х��Qb�L�~E<�au��ߊU99�!95ɪ���a���8��m��V���E��S���� ���I�{�ә���8�>�$���E;h���a�OTYW�ObBMI�\&*��u ���f���\x*]�i�#ր�YV|^��-3�geI�&�?|���'�>�Ǌۮ-E-Cb,�;��]\\��&�S�r9q�[��Y=�:ۊ���Lԧ#g��d,�4X\	8qA�TTY������qMd޻Ȯ��
Z��dyRR��2d°�Ȅ_h?}����c��q¬��A�"g$^i6�
��K'��(��ޑ�)�����|,	�@��kwm)��nP`2233�P{;�ǣ/�C���uH��n���TUUec礈Z��2���yYء��$1?��YL����U����z�V�Dab:�^�#\¹4��be�m���R��@�]��(hF��JD[ʔҕ&�h�ÒQeC�);Q�$�����,�9uD�u�f̃:������� ���w�7oN[�0@l��������H��]sXy)��XZ'�𡶟.�����T��N����J�*��?{H�v8��^�N�"��=��h�>�F<~sk�ʂ-ʞ�/^���ʚ��W.�
~)�|Xgf?,�)���e�8� ��8<!��g��1��̊ �1
%�;�
�xC�U{4��?��Ђo�9�Og���C(NwJ��#Gޅ\dp+��/̜l�-Z ���J�6���a��d�� 3,,��1��5і���o���'�Cv�梠��?����$��Ц#x[���Y@ouT��_���\�R �מW�,ʘ�m�|�Q=�\ҿ�T��$/D���,�u�4��\g;��Q(��)�QjE�K��W���tf�%F���_e���us|�}x�����Xm����W��b��J򠏘�4Xx�ر�_Ѵl$������D�S���Ř�kʴ?,(�\G����i�F�㝌����L�<ʚ��k��dD�u_����Z�%d���c�Eր. �a������ أo�|\ǌ�b��G�Nt6���b����ֿ:ˌ�}��#|ׄ}�L���<ب���t�/� z�i�m�F���~0܈����z-w�\N����T�{ǧg?wN%�1���J-?Q�`�G�N���FK�����7b<�P�M�A������^��\�C객]���*�v &�_[#ʺ��z�����1q�ݻwU��ad�}�+�qX�}�I<EGIA�$u~��װ��&(U�	�<�H<��_�>����3/`	�>Iq���_����3��[3!8���C!�U��#]e	�	UR��U��nD~	q~)��
n{��N l_���u�9�(��x���K��wiM���o a����T�5�+��P��}��	V�-GIk�툫z> �P�z媉�/��%�!�-(�� 0t
�����GQ���O�+4�Ϫ�A�C�a~��몪*E4w���е CE���o�I��!4���:+�� 0�~��d��(c�9�&%ň�-��Z~��1���G�t��m׃��a7�N{8%�5��R*\%�?��+���@�}9�gb61c* �x�*/F�$Q]doŸ6���ǎ
+��̭��:��\��:���^�ԾȐ��U�g_8�
*��:2��AČˎ+I<*��Z�"'��/j�֏���B�2���(n�Zch�|�*��K�x���D�R��#��4M�d�#��kkʄ��b���_`h}cu�� )�߫����sEd1<�W���OAg��v#�Lau����q�?�@Kv���i�-���)��ege��[�U�`������6��<m� vSq��֋oUP$��lK�ϓf���V��Ȓ��#sss���A�[�7��#���/,�ӳ< {_4�������Eʭ1e0V7�[�)]�=�@��rUh�.�:�!�Vy�wK��D�g8����̜3+��-pe����`����� �A����QQFEM$%�`'��<��'���u�D��m�W��}�0�mѐ�����i�ԅ��`�%�W%u�̐~V|B�[f���I`��8��\�h�H�[�:L5=-Pd9 J�=�,���`pʥz8��[�>LV"BO;:NI;�����:!��,u$Z�-C��}���+%JXt� �y��2(��Q�є�h��B�R�1R��須��׮���}�ە���3ێ�I����3 ��� ��Գ�
��<Q:���kx�K�;s�LinhJ�[GJ<xp���쟌�0�a7�Xz 	=B�9�=�픒Č6u����Ð:R�����'"t��[M��
ނ �L��K4�"g�XsΙ�Z0��p�m%�R&)wլ�Os�5c�j�>R&w1.�F$P<��_[S�䟢��yk���>#����~=%7w_��O�ʡ�]y�>F"M���a�T^|�>��8�RH�~5/3++�ִ���uS�$��`��)��1�:�E���?2+l��Șx����3�܀�������bј9��()�߄1�9fD���v !�׹�	C^�n�;4��m��)�����n��t\��1>EdV�����P���=߇!{�G�������.'Ģ�W�t�s!S�Q
����cd{n=�Sy��Ր3��uT���`'����������D�y�_�CJߋ��?��P{�]�*�Py�L�t܅'��@}qR�����Z�i>�r��;c+�G���\2�$a#N�G	���`���9-�y,��/�1��v�'�e�*��
�h`�X)�����</+�����Q����>ϒ��l���g�����!?�n�٧V83� �'���W(~��Z�s�`d�u�A^�
���,>گ>B�Tr$�L+��~)<R�GYp۹AAA�(r��E�j`����?�T1��k��[�Mf�5�3����;��A��.)�ּgfК�P�Y����Ϡ�SYrvY�E��s-6vo���vx�絎6���T7>��^��Z��{&s<�c>��f>�y�PUEE��;��(��xVC��:RhU_P0A��������$⃨G������.�)#.B��:�Q^�l�
��c����9`	��cS�2?e�m*K"������`0�>�?��:��w Eb1f�*<Ƞ%�s*B͖�2�]�09�|���
l[�X�q��}�����^�z�F�t1<H&� i(:�������E��P�4�S����z�f��)N�{q閂�לɵ�.���*�;����J��Sr��0Q'�r�cA�bG VsQG���
����L�#�ŷ=H��2})zC(q��uf��J�ݘ�b���΁.k����J�6+G-�f�e�3y��1*����JD'���uFB�d:*@y����kP�5a���^�\�p:�]�o]�,��ɿH�o��6�#�\���S�6�X�.RS���d�w"1z,�V����k���h�1P� �\F�*k�w�ތ���NK���z�6FG���~,؂���QG;�Ӻ���T���@��Vw�@7����;�7��p�2v�=
���a��ۚ:��������ف�X���e0>���^�da,����u�9���� 7;k���J�x���t�,���sC�M�݃�s�z��ix�Q%rV�&uɹ�r+~�mì/̗<
Qހ�4����r��o� (�H�R�?��񣖆�F�jj��U8C��G�Mq��O��e	�M���G�|�/YL��ŀ�2�)]L�<��2��N�梓x�P����T�B
t%�3s�H��������7b���>p.����*�6�otLcYr�DR���~TT4���2dI->�@w]r�`��n�(Z�斖@�V���RKU�pwI��ӤqBB��ȞF����,<���u=���;K/&��F���~��.ߝ�ؤ���R�*L���8��nd�]���q�1��Τo3L:ۆ�cH9[�ܝ�ױ��"M��:��a�y��<�)yf�������
���3��⏓y����t5>m�6O��� �L�ݧ� `�_�K<Me�#��d��d{��"�����M�w�f����0�����M&*�K~$�[�VdPi�/�c�@�_dh� �2s�u$w�]�w
[g  �:i)���Q9bLGÔ�o��D��9�q��� k8n�x/j(��Gw�:���A���ۋ�,�\]�c�mD�t��o,lP���Tw��0��6���dצr]=]��5S����$Ui�n�w�P���_��H�SO��x���7�%�K�0�V�^�����׫V=_��ę��7�ތd��~%�����"��{|jq�Wl�����ĶA�#]�4�	���(��61M��'O������8�ba1>� ĺ�*t"��Y%A�4|C;�c6�t�����M0��]�!|��v�-xP!0G�eX�i�g�?q���i
}�Li������̪8O�e��A��X��g���Ǟ��F)lݪ����q2�^��l�)06j��r�J�y�s�o`T�1�׳��JSG� ��b��bv>�ϟ&�p5[o`a��L�JF�.l82!3q7J�),��*�}\����y�hzv�0�"!}��Ҡz8����ݷ�p,�KȜ &#c����&\H���0Nr0w���"=�VVw�8i�b@
�m�݉Y�q��X�m*��O�5��VW�o4�F�e��r �+���$=�����
��3��έ���ȥ�Nk9aSSS,3��	��f�Ns�86����Ү�����1�U=���'��rUC����BG{ߙwӓ��s�:�!���%��[�-W��2ʰleUUfUuu�/�@�����! u���܋��L� ���j�Z�P�`�Jy�����ׯ_'U�$�=x��^ۄ�ȟ��.��k��ڙ�;�;5�_JQ�ͳ�4%9��]ۗ����� ,Iwuuu�����(iP}�����"��p�s��eJɞ`$��
�d�bU�3����35��v-�ٲeKe�OY�]�么"���[����j/
��B��5��o"	}YM��A6�rK)BS�P�+s^Փ��S�E(�|��
gy/��g,`��o�1	;�/�a��O[#u:��D��<r{�;�^m+;��?�Ճ����/%�u���о�{G����(�eUT�l�ښq7�j�q�^В���8� ��j0�
�a�0�6�K2q�q8K�����K��)��>(HN�%A��v��)^b�B�[M��,TUPPؙw7�ϯ��cV�iu���4�>�~}�%�D����� ���f�{���>��'�0�:��)�:�25��G��w�.a7�}C(u'w��E�z� �,�z����e���|��G�)/Zt��0��X�>ۆ���W!5�
�$��l�?D�}�M�z��B����T��I���8�'*C�����z�Yb 
u���"c5����s��ˮ5޶\�ޙ�����jqpq��O���G|v��mk�LP�f� s�U �P���;d�0��ka� ��]0���?!?�[p/�ӧ0ȸz���aH(>��m���Ͽ�� �^��0��Uc69���	AE"|16o�Y���d��h���R�^����W] .Q�В�-� _��qP'�E׳(�nI�꧌��e�̲�D��@�B�f) *�b�����������O)�12��󇰨�d��2���T\-�J32��̙�cL8V��q���"C��F�*	����7��t��tC�tVf��M�|�"G�377w�-�G��5����� 8�E8݈(A���x�4i��vڡ��}#7G����Y6�����N`>r�ǎ��\��S�	v���~8���w�(ۅWm,_�N���
h �q�4�/��F���t/�3	e~����[!3"Qҡ�v$U?�i�ֹ���716��:�$�A>R��SC����Ū�5����W�ԙ-}T���o���|�����z[6#dk��O5���"����H��������sĤw�E��oC���I�;|�5̷��ѧ�ڳ��M��k��yI ����T@y���K�c3}}}��U�䩅�<�ga���Ls���Qg;+++��r��8_��pX�~=u�л�D��C�XX�w9bd����.A��F�ڰg����`�sc-Θ_--�6�:�e���^;������r,��>��y�����VB��y�LC}���x�eGG��1&��Rv��i�7���x��;����?�,�W*�FG�Y���l��y�
�1��;>�8zX�)��$�{7�L!%O�J�s�ςjbz��{	ƫ��)��d�oI;���,���N�5��BAp����\�+�:��:VB���D�,i߭�3�ԑ�gϞ]�:�Va�Sz�1$v�"_&B�kXs��I�|��h��=�`�Z�o(�VGO�z�q	�OKZ������o�������:9��,�%z�;���ob��3� �Cǲ]x�"��d�Zd���}(xE���:��ͣ��;J@�}�$S1����9s]z�z:3��A�7]i��Y�3;̉5I�X���tP���#�Ģ�I�MzP����W��R��AR�333����L��������x$�*�� ��^�Պ)�O�w��Y�����`!����^ŧA�姡��F~�+���M� �����?�c���CJ�W��h9@�7����������d�c��@x'���~��u@�E�M���ɫ�_Q�-��Um�4�!�Z����\�^���؍�r�@"���ȃE����[X���%2�z0��-�}d�8f㎸\ޠ�~�a�)Z�(��,|��07B�0��X�_��1�
`ǟ�J���;A�<M�>���;���=�+u�/l*��l���	۲B�<�������S_��	|���^?66vU�� dD~����Uw:H�w�?��b$7�4�[`t|�͝P���U�7o6�`l���=@�7��*�~#'�lG �Ӏ��VO^A�3��>$A��L v�sF���YFՐ;�O�ܡS�����ɨQ�üN����Q!�y����kZI���	�i��.�/�0�ȋֹy��8\�UQq�I9�:��:�
�b3C^�#�=v��E���mca�R���m�9���[��*����c��K��JKK31�g�������t͑g��H�> uX���<h)�ؐ��d�z��aB��7{7��M��A>C�xz���f���Qбj��hx�<�W�_dh��?Y�}R6��6�{ hh�W��, q[�㗜5�To�z�� t� ��M�	��Ѧt ����3�:RpP�����}=>L��N�- �{QR�9*K�����3J1���0VOޅbD{U76�8p`2v��B�7�N��?}��2u�:4�����ZvVm��V��oA6h�w<��uv�%�N�<ٶ�T��K^Nt�q����,%�+Թ�U��3�$W�%0����!{�@]�f J�R0v��*///'Ї��8���F���6$�=0:�+\ɞ��ѐg���A>��	7W�JK��h����	����L7X��3�L�g;�O7����q@+���wyV�ú�t��@,)>�������H�򧢼��uK���`a�ϧ?��D?؜�ρ]@̛�v������c!��Y�3�<�\f��.� ��o�# Cμ��dx�����㉊��U�j7�pQ3]�\� d��u��"�XvTvȹO��H�$a��!���ܺ�7��eCrT�"cc�5Z�*�"�$F7.����ʠI��,0i:�6"��������r��B���S �::�i5/Շ���6����(�D�T�U������ZdǇqCCC��	��_��?�w�)�{�Z�J~hʁV����6z۶kjhL?LuC�PZ��`�L���)�DUP���!# ��h�>��V�wf�`@󥺄�����:�a�\s)q��dBF~����X�R=LDpx�����L�����6���o�ԑ1o�Q���6��6��S|3�B�j�?(U��1���|�#G޽���DCf�mY�o1?T��4�Y�r���g��� ��Y
�����8h�����Ti�I�x�u�!�&�e�����.�V��a)}of�8 �΄�*'	ŗƌ�s�C�iK�J����r��!g�g����,~�Niu$�r�u٫���c��-� �y##CL����i}�DYHd2��v�� �^ja���9���\ZQ�Lڷ�i;4�<F�Г �q9�����0~�e�gj���A}.�ǙZ��V��ToW��� �O&߯�~׼�1����v-%?�tN�Bۉr��f����D;#L�(�#uO�K�'��i�6��)�K��<�8�cf�;2���-̱4�1�+HQ���n`�9�Ȅ)�oZ�} 7*�qG�s(��7��&)������GR$�����������O���>���w��r���6��i���u���JB��ώ$d��ǀ�����Ԁ����PRn�In?)*�E��	��p���=�x�5	�Av� ��/h]���c(U|X�aw�r�4�O�,+q�&�wy�S�s`N�&���e� �ƺΑJz2�y)L2)[��n�6@���*kj�O�4in��=Bv�-$���F	��� Y�8��Z4�n�m@5�̡�H+���	�ԓ����n�L�t��[�i)��e�ھ{�޳�����h��t�Q=�EG��U(�ZXx�5pT�-�����m۶堺�Y�<�u�݉5��!�Є+��O��A�E�]�'����X�x�aH����^ۏ�k�;5�jd�1r��w�Z�MO@CZȚ���P<љ�y���+��h�V��. �%�[�I�5�DQC�ײd��&���z�A#�	�K.�#���3Ϟ<y�vp�;I�R�q��,����D�[�y�:it�՞d�c�b�uf߃��(�򤚢��n�Tt�#u����b�����%r�
w_X���w�2r�F�ҫ8��5Eb����ڲ!3#������70�ؘ��{I�*h��Uy�ŸzrL1���yTsȣn��>��ֽ�Ej"^���p����vD�K��a�\gcB����YWt$�ğ2���gd�l<�,��jg>�?`$u�V��c��ܒ�V���,����9S����f����h`�`��Q���ͩ��)��<0�܂�Ў�=ʱ�Y�usW�^M�+]ۊpF6�nM:�ҍI&�Y�Y-���к���u�%�Gl� v?ǎ��-}�������D�mп�������)�$�g��>k�=M�ํm���dD�Ni{,���.�;@����x ��%�u� L��
��|>a���%���@=�Gy0���ݢ��]�ϸ�)������	4��!�-��8�ˌ	M�3<�Sr$�{�,YX�j�|�Jo���(��Ͽ��4JH�|���E]�<��8;�Kt'����e�WѯH�;;��$���|(Z �8���H���r���{,G��2D��tu�v�r��e��,u��� ��0ژ*��Sv�Pt���l�2sKصI�&�;��n����$ Ey�;3��|	J�1d�����&�o�]��(t��TQ/FO�n��f���_�
�ԙq�>r�l*3��B=�Dia�|{J�$�����Pj�BKآJX����=�J�}��CY�=�Z�ZE���3��뙙q��^Z'�<�ɚ����vm&W>��	�<ˡR�Pȿ�*����ɕt���݌���a�XǌIn�W+B������ఈ7|<��4R$�I����of� N�B��vV�B;*���&w�4��uf� ̿M����RR��0����u��=h-�C��C Æ�'K�T�BB��&�j"Nn�=�N�L���T������mu�֠q`�8k ��-���)�q���8mI��`f��r�г��������u^��[L/������F��RFF�u����9T<Wj����"D�>Y�d;�����S�2�y�S��KF�
�Hw$c�b*��Nh��2�r;��gz֡�ȃ��>ة���g[�h���@B�")�0MC�����zw+`���B�!ؐ�'%O��g�#ϑ���@'�s~�k�F�`,?O�l(`'��_�R���r��ݷ�E?Q/'}*M#��慰Z��{r�q�w��^��9�c��R0}��4 o�P�:Z$�y�1a -��1����+v@RdP����xĩ�,#�C���w?��82�w	�����n�d�|�����T��S�d$EB����y�f\�+��|a�^{��Q
'�{Ӭa�jZ8b�c���3{7$�]B� �Z��]/37��d�23�gg���1��sR�@t��T�5D;�u�dNJ�ϻ^5+����u�y���.,�L�"[� ��B�<Cܨ̾�Y]�<-D\6ɼzXX��km#:�ƍ���vn�>r/~ރ�Sd��Zm�x?�s�l3���d(�6(�Q:p,ی���e�/,!��l"ET�&���϶�
{�J1d8�oñ�d�\�9Z���q����$ _ħ��w��}�����U��"���W@�Ői�0L��!�Ts�t�^���PCN��ɑ�E��A^^ֽ{�W#�Tj�Ni�����-�Gӫ: �H*,�\,
�tm|Lʭ�����H�WF�A�n|C�l �	<sn�ؘ&�d(B�K��؝��fLu�K�f!BAkԩрtD��<�����f�+���r��nZ^��R�@�n�NLYN����ت�����>��h\X�����E\���?B�JI:/P����>%�K��9��ƪ&G跼�ϴ���.���g��7��n߼J�F��ʯ�j�?���U�%��/���~o�����ħm���V��vm����k���S��Ǎ�iI��S�n�3��������} ���/Z�(�ǧM~�+��B�/YQ[ŌQm��0��r�|���Eb酐����D��4|<:{�A���62O�N��n�rwj�\�cj�+>�KKP���;�y-G�'6�z�i�D!Z��X���=���K4R�A`|��GJ�OL��:khh�U���y)��H��ce���d 5��_��@�rI��� �Ϛ�t���D��O�}����&�.�I<� B���~�H�~wn?#����������bb�ҫպ�ۑ��a�(��z�� {���5��Y /���Gs�� ��!�ai�W����w�UD+�_?ņ_Q1N���"/�MV�x4����s8�v�A����2c���rs���3�Ô��wa%s���N� ~f1_;��������)�C���b7]xE�'�S�-����M?�Iou|���[��W����]r!P&�4��$-��n\�(�����~~�߭��jL>����k��j�Sz"���X�u�4���	ݯ ����W�:/@i4��d�PB��ĉ,S�6������r���s� Ȭ ,j�i*%���d���6?S}�i3/�Y�+�\�3H�<���c�^i��V�imZ�#��	y;���t|��c���,$���uw�H��;��s�u#�K��ў�h7}�W�wHZ�6����Z�(|`M	�<h�豈�F�>%;�^��/�?a�o�9�wEj� �&n�,��~�h���q��u᧟��s�U}m�R�V�-���H�0�{�u& g�nbjz��3����d����s�a����:��X����R��/���w���v80���9�)�Ȩe?nf�����H+��X�bV�l��$W��I��Ͻ��pY��=Ym���!�.�0j\�'��f�������p٪��U�5���^=gq������T�ﾁ�����+5&�R(���0�*T���@TΘ�p[�	�=G�/�8?��j���~�=͊>�kw]��M�u�L չ50gw�4�8���C�e��j��i�̘�ͳ��y#��,�ԇ�`>W�q�9q�R_���>ρ9u03��7���wã̘���VR�>��WYW�ԕ��CG��BS��B'Z�� A\�������Qv���T�%�*i�eu	j1�b�F�Pq�@A���(� ��u�	�>p��}��ܳ|�;��{�O�X�P?��t�I�a{�Q�~?c���;�ˊ)��ɍćtV;�.��f����^���:K�t�����B����~d~ӷ8WB����ΡdH`�]����P�+C���qYwMdz@djw|0��6t�իW��c��0���R��G��FP���oM��mf �EY��$�Ō�Kc��Ż���9���ݓ�b�?|�Q
�_��V�:PRb�pH�ڧ4���2G�}*��2����g�������V�4�[ ����T"�n��F�C�36C��� ����ս��k"��-L 3H@8�/�s'S�X�]�"!���_�	Y`�_MW�,���\<�F��cnl!��ʣ;k�GD!��s'�ȑ#.�`���� ��R�=^�`l��~��P=�}߄J4v�\��y�b�Z4��D��0`��o�gI���;gŻעmR�F�;��N����JJ��ΎY!�e8I��è�ą���w��G9�V��_�ݶ���Ũ+��]�e)v������V!�=�n(<�R�#��h}��Դ��䌞�wI���$;���L�:d�<i#Sa,VnaϺm�H��=�a��T{}#�(r~��oo�| ���0;�����k�M%H:R ����GB3��Z����8��Q[�X�W�mh��%1Ke���q����;�.<y�u+ڐ���o����=x�4����.�p)�R�xW�����C6p���uO>[�Z<k�c���#G?�o�o�D��;�*��c�I��_xR��sF"Y�v�4����{�>�! �-_i ���˪�B�4�R�5�M��k�e���Q6�.���0-G._~T4v~�W!���m	R:�)�r�n���������CXMҏ2O����G�pj��V�Z��b�]��`4-����?b��]���Dtj�P�<2]��U�-���;gb�Gr��(����W�n,B�bKr5&=�y6����I��#l]q����R��Z(���-z����	��� ��{��LUe�f`kB����O�)S�*�x?���R�NEW)���^�♼N���ܯN�v�Z���S�f��.b� �j�Z�܏��<�%���r��`ΰh��yUأ��eꖑ\( �u�]q�E�@�h�kj�9��41K>	�n���Ӎ�ƣ,)[�����^�_s�j��`'"@�Wmp�]��b�
(X6z�����՞]?�A�0S�`$|���Vnܛ��8$�I�S����\]�O:1���!�C�7U��/w�+	δX ��Kt��ء
��J}$��!���B��k�bF��q1�UEEE�h 3iN����JM�Ʌ/�2l0��r���FVW�k��L���Qq��l�n<�qCG �7ۡ��?-..��r�g^�u�Ɣ|:O��HP,^����~���P�>Z˛~��JQ(6��4����>�?���zo1��O[���t���$	V̉��e�a��i:�U�� RX��J���ܻ����5�*����pLB)D3k�i��ZV�ד�COq݄nU�Q��Z�x��m�i�,�Aޑl��.��[/�r+�j�|����p-k�y� "Bݑ�a``��V7�E�;(�<|����
�jl�@N �u�Z��@�u���`��s@�by�y@Kl�b��OԿ�ܶ��r��l��'�(+��O��GM�%���9���-j1����0�������Q��2{���Y��n���3� ��Q��.����yyZmc�tҫ��wbO-�A��"�kӚ
�9�+���&�����}��a}�@����4�zTep�fT�<��ď�w�ܳiS#�9lQ�p�|3�*��#7!�n���0�s4�4Å���y�T���qu!hߔ��Lk�}���ǅ�^UՙS(���^���|�x7��U��Wr��|A��(�B������ၞSvEy�ט��S�?���ux�!�-��GW�^$A<�&�Xxy��XKol�A��T��!rFh�y�k�:N���o.�@��1E�����Y0R��H52e��S� Ъ��xҟc�qM4���-L=�%AM^<d������������l�T�hg�i��'�H�	^j�{&�^@/do�܀ :�t�Pg��2 �6#�%�+�Z�s?gDa�����y~�F}���OA���� ~�ԠǷ��J�ہ��]8��k�������u�����+�1�Y��d�����'N�]�]�7։��!������G&L.��!ЬA�b7�s�^/�x��Q�,��"�pߛ8C,�e3����>��kf��FcT�ݾQ��Zz3j��b�z��jv�J�z�)��W%P/Z�*i�iq�
N I�C��k�����7
BS�R	Pc�j�ׅ��""��8e-0�� ���)� ���)�u��eHr�g	ԣ��z{>s��t��\���H�	O`��xbe[֘��x�k��N�x����*v-뽠��n$B4�=�[|��va����y�S7b�V�&98b��%��ɏԻAU�k��m����<�p�A��}&�L�8�[ox�>'���T�]�����V���Mn;R��q�����`(!,է�B7��i�h6d.���/���ؙ\�������*k�0�߄�Q����_�
���)��Ho������Z1���Pp}8�W�ye��Oڄ�2�t�@�Bڧ�rYf�ծ��a�G��B?�8���ě�eL����?��F��#A=�m�	�B"���)�"��=�,B;NXd0���S�m�GO�K�����,o�`Z��s�w��8ԖG￨�y�5R�&Hx�-ۮH559���>����xJ��e�Uea��+�Yꢏ��-�q��������w���=�Y	L�,Њ�4�wG�n�Κ��\5KJJ�I�!d�3�� ��0�{����< %�UC��ȫj$]5�L4h��:K�'��sR!���\�@��ڙ �
�����'v�d���:ko��a5/ca����!I��X6d ��Ȟ)ɼˋ������
Y=�44����/�d��u=����v$����.�j%*�f��%��1g���Bt!��!�UOzw�Z�V^��y���'�v+-t�W�9�[�qԞ�H��~>Ϻ|��KAJ�${}K�cW$?
vt7��a��t<J◑�����Ҕ�2�=�����iҸ���~u����&8�*���yT���N�D*ډ��L���;�F��	|5}�c�!�b�8���&CL���	o�~Pc߯*��/��`�PGn@��I-�ɂr�m�]Qs3R/�n�� ��qM�k>��ء�e���%I/�L�O��iX_[�GkP������K3��Ł�Z7A'nW�Go�ɼq�ShvuԠ���Ҳ�>͏
��e������Sw��� ��|����C*l{�I�FvN[���h<�2'�Qn��-���u-P�c�����]=4�	��T�'<X�Q5a�R��D,@D��t������=_pI6�����l�"q�t�g.(Y������$e���x���p� Z�ftҲ�k{�g(��}��U��gzk֭.�kۢX�0�5}���bh-���݅�����jz�^��|/�vز�|�o���Ƒ������ PK   ��rZ A��?5 �J /   images/e0d6f4e0-adc9-461d-95f3-67e9d6b55837.pngT{PU]�6��GZJA@ �(-"����tw�#*� ��-�twww�k��{g~fBX��k�����,>�}|y9��((�k((��`���>eT ����iأ��$B�P���R:H�;�Z;8���8;;�M����m���v&q;"�QP��K={��5�����L��n�z0I��}m"ii�����ExOx&��_�� ������hSO����
��(M7��ߣ�Q�H��=$�������[��ܹ�\%q��L���O<�c�Ċ����>G��@���s� �KG"3��	���^��
!��U���i�=�6o����E����D{��ܴw6��bݕ�2�a�����e�p`�p�/(\oz߽{p_XE�$�!`o�@��ȱ��HN�"�75�
�y}�ۃȍ]))��W>pzz��������dȦ8Ȍj��7C�����O���JVv�P�ob�N�I`0[v�5���Ϩ��ug!��k}��UI9��ddJ�spd���������}��-	)��۷�����8��\���R��5~���+[���$://�e<߹9��˳3�9:�q111L���e�L��Bu6���@�?777g����}B��Y���1�e���v�.�kS�$R..M[Jj�:���h�j�ʡ��ӈ/..���������*X��
��qAFJz=���q�+-�m��,'w��Ç�����������^�""�{{6 �kCّ��(,ял��n>�<h�!$��L_>�#-�J,�ƌ�a����V˟'p,����eQ\R������%Y�@>/((���%kddd.Z.y����QX�I��p�|���{���8%5�ȼW6JE;�� "�v#����:$��/�;$J��М�Z�>����橱����EF�^��Sn�6$��S?��fag�@C%%�~�$<<���F������3E��r���&�ֺ���W����Q9z���$BG����V�ҩS�P)��34|C>uy�k��9N����:��F�Ǳo��sqq�vt�C���ݸ[X����w�i�m�d-���T.���=K�>b�R�o���I$�)'K�������yyBo6<�����eB�+RG\H�'��I�Ҋo��w��2ڢ��I���%M-����Ã�;�X��v������̞dgg�m�d`d�RZ��u��O:?������۟�wn�%���ӝ�(cA]+�)��ÃKe�>Hdi4ԓ�o������p޹cхMBFVl>
��*/�oV}���w�G߶�/A�>�~�%ݟ(�>Y���d��K�^Q!��I��($�7?�r�B��辜���]�KKK�N[c�^�ᰰ��ed�IiMă��8�U�ƛ���C���5~(*]28���<G���I�?��
�u7��O�"�.��ہ�_Dd�����ί����I�Ʌy��؃ֺǛ��!��^Gøttt�����wqs�y�21�`�|�0��r���-E�h�%>V!3�-/��j������.O����2������֮��	__��~�T֟k�a�1��ۢ���^HV(�Z�D��Bس��?W���EK4�,--�5V��2���~T��b���W=wI@)��������_�	�Ll���5J�O�yF[A�۷�)S}P��PpK�u��D���0bE����+ Aع�t�������d���u��p��?11q�7*��i�<�@��� ��μ��P
�ܟngOL�Ia��נĎ�d���P`~�w�tu�q���\l�((���fy���b��%�s�O�ӄ) 9A;��;5M8�pO���@@_B���N�<c%�}��ξ<��0�xi1Q��t��}pp�b=[�NUI�K�/6����y�>oy1/�Lg?��J�meJ����e�˳��j�:���yO��K��ض�*3i��Q���p�/��ι�x�y�ssz�V�!]O���������8���+��¸��hw'D1-��=bb����T|�44�#~�/�~[�2�$꣰�B�&h���|���PO������
�=�����ǚ�>�<�d�22X��������GČ����,�������J�_����J��$1��Xv,����vT}E�`@��bi!9ϸ�Te�н�k!�::T�}_���hI8[����nJ1�a�s�9"&��\�$ l�W�]po����x�Xf5cb��i{B�����\�Õ޵�rd�T�N��`�M+�d�ޟ��zi�դ���p}�4�F}�*��9B�gk({�M�w47?1�׊���6����VE
f��\R�RąS�p>޾�!=}J���S`ўXa7/����b�=��e��ܷ!&F��B��^���5y��A62%�sC?B�>$�A`�r1�ƈ+	%	�}B�+��Eho�Jm}�x�(u�7+&ǫYg�Bv�/C����eH`�gg.2!�]��2O��W�b'}�d��PƶR��M���Wދ�o�v�����G�'RV�����bozzvY��|���c?���Pe�iU�s"�[t�j�d��%�Kk�P�F-��j��HII11/đ�j���Џ2��L1QQQ�hE�UV���prf�Lri �8{���XA,b��g��d���c'�
�,�V��^�i��<;+��T3�?<4X�����K�ɴG�E����#��y �T��X2�+�Ȼ�����o߼)t;6���`���6s�FywFiE®���g{�g��#e8�_��7��l5z(-5A%a��o"�5�J;��g�j5J�K�k�1W�*"��u=M$�J��`�����Hnj ����}@�P�]�S��2���$�r�w{_�!4M��Ǡ%�?.��[B���/�/q(ʉ��L۩�3��h�)���1�xGL&�iT.h�����M'���9����&����6 n۫c ��`�a�h���jm��D��O��$ٳ�Rur����n�і��V�2)<X�l��	#ײA�"ؑ�eI���C�ʀ��A�p9�FR���;j��j��`T�ڛv�Uy��N�@1�����K]]�斖�ؙi}��ů��W��77���c�M捷޾p\���:n�C���8<��Ch�ի-X���?%JX�ӌ �չ�������K��w.;�F�Ɔ�$ɓ/���w�ɗ�ҹ-I��[�p'%н��zC~��� ��Pts�6�*W�������;�����T�T�+�;��$�%YY�`z��W�UY�5�F� ���VJ�9!�B�l�Aݝg�#ɣ��w���\I ր�>��+����ݻ/��Wb�7�p����`v�?Y`M
�H�k��Kjs�~B�FF� ���&I11��;���S�=sp�bL3i�;:�^���椢���W=��j�N��Z1йJ?A'N��U��"^yjM�x4����λ:vvv�;���/���k�\8`����u��B6�� � �9'^�9-������;�4���.\`��6��u�'���e��P٫989� ���{�5$d�.|.��ݟ2�Q���F~��Yq,jd)%�ټ;˧�[��7
�[����PA{ׅ�âJ&�!��}���T������#���,��,�*���e4�ť�}�L�U���m��~��z�%�*�+1L�5`J�������R�;RQ���q�_}���b���$"�N乺��T�Ķʼh�,�ˍt^��}}+��b�-_�"��v/��_�U���+ F!��ǧ�9����ר�'>H�#�#�z���,|�߸Pe�88s�	����Ť+�8�{i@}��&��y?==�����g�O��	a��%�lA\�����5׭��6�4�|L�F��дp�[>zJ}��D�ځ��t�s�X����e�/6��id������Վ-���w�'ı3v��f=~mޓ�ҌD`�)7wK3~�I�%.��/vt*�� �A�9��i���2u6�~�
u6%�ћ/���mѬ��Y��^�tţ�G_U'\<$� ��B��~�ܗ@�����;Հ߭?��z�K�k܃�; �ߚ� ���Yp��� HJ��v��&5\o[�S����;�4-᳉`�U$"l@-�~w3X���G����ܭ�M�
��y�����M��Y�w�^���k&yᙍf+'��D*	e'Ý�`X�h�ZqJRBO�H⠛��gU0Ԙ�B:��̣0���T�(�P���%�n�_�-�8CCG/�xl�$���;Eߟx�G���2�_	B��Z_�Rǒלu#�a̂���v��z�/�@<Q��vs�P��4�m W��i: �]W8��j����l��-��ޝ'Cҭ�P(��Z�8cݾT��ެ=�0�QŜ�Db�nUT�:Kv��ӓı#�gP��H�����pCA��	�,���b,�������ܺ�YXx������۷���gD����̹G�n�WZJ�se׀�ߊ�ٳg��稾��8�L��'/�A��9])(Tn���%c��;��X��N2�=C]__W�I�	����|��K�d`�۵�CXj����fG��
�ly`�&`˝E���y8?�~�,K��zU�Bwo�i�e��+�~�j���4����A�-�w�ׇ�U%���8q�W>�(AԕjK�D�f�U�.�P�*�w(�i�Be�j�9�|��������򉀮X5M�jjd|q��� ͹>��P3f+�U^�Y����|��u�B�M�RjB �����Bnl_V�r���~�����6nZ0�1������W�^�!����+�������N�U�ߝ�ei��J��9XXvm��8��>��x�q����{O�+3�[�C�+ſ5�����<���M�2���������|\߾}���I��9~˃'O �����5�?~���_�+7��P��w�tr��$�{><������]�R��F�YL_(���b�i�o-.~JƦ��޺!�w��n��p}BCݽk;33���~��r|cs��zƣ�֖,�@�PP �p�	���R�̯����ԶY*��������n~�)��a��Dd)*��5ZFOaSs�蕌�NvY~b�H�	�nMל"SN?b``�����ӹ�2Yl����w�/r�G�y�yw[�UJ����6��R��E`4��GNA}u2�iz��;լM�
$u���I��<���.ZE�T%[�.�tJ�6
ڄӬ {�/p���C����)���9yy����#
,Q��V�^�	>;{��ˮ�L�����nxCP��M4P4�Q�\�>�O9��)tH�ީFU�E�J4T;�$,wGn�[ϊ�K��3�EE�8���ঝ���k�Ъ�������\\�ΰ��~�(6�e�(�([^ɣ��\��Gܜ�_��di$�TQ�|E�C.���@�͗�V�D�J�������^khh F��?=�1��X"�}{t�P\R���� h)YY�c�X�:7��@X)���6��Ɂ��@�WV�����h�����l��5�(��Q#O���*,L��0�W�^����N�[�Z�����"gNt��_�K����`�R*���1��=�I�RS�|�uM���u.�q	#�uOW��=\D"+�)) @��<�ag*�����|4�����W6R! ?�7�Z5�C�?���&��G\�$k`�)�463H\jeq��=>`�>�����\Z��y��`�u�')��k>* s/�wsppT;m���kkz�ř�~��]�Ls����U_���\ZZ��۷�������<hL��8<=]����� �{�!޿I�W�E&��27�ԺD9�V���w����ڣ�m'fm,{歈�h������UY�!���ya=U��k@ "�����m���_�n��|������3�����[�0Y��~�G�t��A��Y�ϟ�'��mܕ22b&ļ��8Aȑ��CT�V�v` �s@�[�z�O�ylL����.�Y'a���Y^���*���� h"�S=Nt��̡�77�C���̤)��RRS�?z���U��B��_-��5M�I-����P��]~YH�9~f����n|�mͻ�הL��ᯖ�>�/H � G�P���<�&���u=.{�Q����M[��(`3��>����V"R����<h�����w77,,؀��J7�� %҄I�i���n_���pP��@��]S|�*i,�~��-�f)2J�+�m�~����N�|+��G�ݻ7�$i���Y/����o�W���SW�qUW�T��u���襂ƕcU�?�����
3$Z����ao��*�~,�H��Pʹ�O]�!!��X}ro�f�ilZz��e�j'H������CiE��V�D{.���k������;˒�t�b��\��3Τ����h�HOo��뮮���A�JcQgP�;�~:1�w����g��������������O{�h�؎Հ��,%Ʒ1SD
R�>�ʳu�XM���\���^�L���"��֠����U��]΂�FV@����`yU���f�&��ρ9R��i����\z��~_�`ZF�Еb��D+��Vt/O��_��U1^�(�a�>?F#�Ł�2Z#�07g%��BC{λ��.�h�:��:��x� l�V��G ���=E���(�^8n�{":��X0<s�M3]>�5�s#Z��g�^^(�=x�S�*����=zg{����d+(���L���Pع����Ϊ����En�c����,&�;�Vq���������dd�q�|�=�_t]O���d	KH���(qY���ק���a}�-���	
��)��.�"�*��w �<�!���Dۡ�1����2�V'B��0��o&�l9�^�I,ʴ'C 4q�_��@/SS�^+c
,��>�����ߣ�;-+���R�3?z��Vԭ�P�v���[�
�I9q�nX�ږ�$� ��ժiIeyh�g=�S۱Rd�O{�0�oO��s�@O(�G�%%���枝���Z4x{���'���Ӳ}��$�/zJ}:�L���H0�DT�մ�g��ߍ�
�݄.y�7��Q��}��������j�ܕ��Y��˗ڋ�6��F#s,i���zOa##���}���z����ű��)~��n��b�A߷���`��Nн�{��<6G�98
V��c�)�\�Lqm477o�ޠ�Ry'X!��_��/h���7��%��~i��chP��#1 
M  �����eR���������i+f^��WWWƻ��9��Q���!�e��9v���*o�,����?Z��Tъp�D�RB���d�Vq���%[���YKe)-���
�F���n�edfvNɎ���}���s��,h���v���kp0#���%C����A�bCyI��� ��LJ��94����@�U_�k�R�q
4���^>6_��ȡT4��koa�s�=ƺ�Yr;��������J���$^�G'n��~�$�@2A��	����u�x���U���g�AD*���(ĽD��w�_(��F���e�6ܶ@?��`���ג~���J�vh��d���3[>k�?��?�N���B����b���^����a�&�%�>/���pC)�/���|eFz ���hE�T�5�-�]o��vjv�9�KL����3�$OON���	���<<=�Am���$�VL+.>�{���p��1[�f*�v1'9t�  �3����Y��	#�v�IJJ�l����]l���Q����ڕ�^�kc1_�,��H>?^�DRu��
��yYZ&Fƶ�ERRi�kD g�EH}��ѣ����<y�zR���i`���/�rs-�,��^_��oe��X �a<�&O-`Ә|C����%%%%>�Ƕ����	z	%��ĵ�)��L�:=<���;�&�UZ���Ǻ�<D	4�S�+"��X�����x񢳷W��'QPt���$\xe�ݻ�}ɒ���qg@���C��jמ	�����(�ߥكw��rݳ�x�	~�O_H-EC<ZM9k2�Ԕ�jDx�<T �����8��v*ώ����naY��cf��?����k2(lڒAw��Ng�Ł�p�V��FY���1^^Кi<�.5Ғ��lA���B\\H�i�ٗ�đ45����N4�n�M�w�OO3Anh�Z8�����)���{Ine�o�.�AG�ԣ���3��7�-G���ׯ_Gz��C@�2��lt�5���r����*�i����?��J<(��C	����!L�{?^(��3=λT���݂[����p����(�t)A���5�i5U��3��b�6�+���vQl���p@����c��Fu��o��/8~sE���]�����k�G�lBd����ņ���P^^^1F��������v< v��������|�)��rU���v��+?���u����-���F�������8��c3%�e$3W�T��3�N��r�N2k�y�8�:��fT�7@!�q4�fT}�j$��*�Π��z��]#\qI+��r!#���t�#{udF�������f�U�:�#�ֽ�������XC��8�4B���")�:)��Ss�s�ݙ�㵵��V�/JqU�և�(tqLLL�Y��;�ӥ�i��*iO�*嘃�u��'n�RE���J��=�˄K__ML���
KJ8���p����p�g=%�[Sfdll�r�dҺbM����Ç"<݀P�jqq�~�P�U�uֆ_$5����\P��4��;k���V�x�?�HP^���0ؾ�����C��M�~H���:���~���m?n���j$_[��*_�t|�	h�����Qr��l�d��H���x���4[��&�~���p�p2�t�is�#7��jͨ����<oo��xv�MN�����ݲ����kP�!��pŕ��G� g��I���y�KHR�����
jhhxoB�5]զ@=��w�Y;E<��]_ko�
LS_�6�4#xӒ�Y"�a��:�kG�$ ���ޞ�PUQ��������x4Fĵ7�J���E} ����ED�++ ?Ň�p��s:m�gL����9	Rha{�g|��2���`��*��M�7�;&�?ح��ɜ�����В�`��3x�=9�}tvW�Sf� �� z&&,�T�t������K�3���>�
�;S�:��(^U�r���;�4$���@W9�beP`�ŭ�~������-j�W����4W���=wp����ݝsN� ����T�r��c�|����z��(��rE��g���e����`���*�����Ɋ���\�K�������A%�^��)f~�(YZ���:.�9�)��0���O�X
ׇ����6����Y�+�+[�9����7�~���,xV���F�d;�9/j��|-���edDDE�6 xR�Uo캕b���VO��Zj����m����-�N�����@�{�e��䊉-���3"H��7YTLth&C|�]�0q]V�M�!�/e^1�vvOA/�<�%$\F�po�	�b�ks$Ϡ=��(UP �#s�w�o���3ewȮ͙|���"�e�Nȸ�5���t]ިo����t���T ��@-���5e�PX���C���$��aÉq[ ����Div۩��?1����>�K��k�k�]L
-B6;�0B@�i��N;s���'+�*�Ip�<�u6��4$�ߝ�4c����F ��+1`G� B��?�M����8[="'&n18�]l%VΝ��9�7�D�#�H�Ҳ�׮�V�gy`�
ϖ ���U�������(�Q+�����S��o�Sb~�yx|����
��J�*�y��`SW3�I]��Z�?M[���˕���1;�rxU���;�*�H$�͛7Pm�W������ j��. M�Õ���դ���Z�S'P�@W̯���9���5�Ƹ�*���m������)� ]�H�§?w�z;[J��=��Ix�"���gC-�;+ف뫫�9_�ʣ�o=���.:��Q]D�\���x� D�ľmLo���ܝi[�G�U8����dR��YQ!�t���V��
1�c"����� P�^��8�Ò� �k/wj�(�������<�~_۔�� ؋�ѣV���N��w���UK��Ltz�X?[���D@�t�?�ks��&g����H�I��J;$7H�ze��(��~�H�L��ue�@��AEG��\�30|u^g����0�n�d�]�no�(L�-7�xU����� B��in��c	��؄mc
,e�c�L%G���F%�.���U (��gb���n'[�%��b熉.Ww�ě|t�4�nʺ?!+�G�������=a�E�_��j�Ut���C�������ɓfc��|�����?��S��8$vuw>�Ų�������;4�Ԕ���#�����&_���x��.����*�|q�d3���mvs�de0l��ѓ{i����UoE��Π�������Oh��<�P���'�V4z����+�QX67���>d_,Ο���6 ,K0)�t�S�I��+�V�(������o3+{�[�
ܱm'~���Է�:�_l�,f=Oi@�\�+#�T��G������ڗp��A7MC�+��N��m�EG��4�+9��L��$�	�=�k�P�����4��j䨒��9���8k*�a߿�}�VU/3�~���\N�<+���b%^d-����Z�}- �R�1���RS#���ߥ�����,���4P�xtb񍍍+��2�G)��i4@&l�ŏ�%��6�<�6��i�@��3�JI���Yߦ�߻�l��n���L����!s,�#(�����
}��.{~��[�����mЋ�������ֈ9�D0{0	�p�?����'̙ix`��[e�XTT�w��Sz}��L�ߌ�3��'܂���{dd+�c ���9��	�j�_?W|�y�����Z4�)�'.W����&�z�2oZ��<���'��������Q Ŋ��h�Mck���G�	�3.���VX����?���'�<��h�^�����"�槂;Qh�jcv~zzzO�5�a�l"�չ���8��X�tS�b��##�Ք�������r�@W<jkOg3��o��5v����wxp�́�`��flU�8R7K5��А����*�ͫӝiP���Ϟ�"λuՋ>|	|]��yyb��;��{���aҟ(
�1ٞ(S��	?::��E���^S5x�D�4��.��U���&SdD��aR
!YgddԲi�9���Vv~����`}qqq�p�Έ�Hmʹ��L���\݆z+{�^1b���5��XN��z|6gA���񮡽-�%U\��O\�y䕔2~�<7�Z�]��J"7r�q<���0�L�_>���L�����(P/��m�t�MKlS��;y>r�@*Y�3Y���=�蹣1�J��~�CY���6� ��i~�N�iI;���j6����>n��޽�3u��5����JK#�D�����1�hݗY� R��:R9��<�����x#����+�h�/����|��~ �7u�dekhO;mk�	��;�޹�S9I��b���|��i���sӬw�3�>ѓ?�yk>]����bbb�lWi����"@T��o�Ԋ�O�^((�l����I���ߞ���:��z�cF�z	���p�r�bH���tׯ��ɨ�$����Z(i�vq��S[6��zXJ�U�\�����/d��) ��������nf��]<t���b��`��T�I)^��۷����ᜨ��Yi�����?ֳս�6�¦t})M9�j�j�h64�[CeEťD��W ���D2�"�����c�Q4��[i��U_>�ʮUf���[#X�OD� �Ur�2
�N ��
���*﩯pҳ���)�ɧȠ噘��::;�ͤ1	���JxK�'##���̤b����%%���j�*f��Vb�WQ�<�K֥����Ԅ7��c������>��,�痏�W��*�D�i_�������zy݄M��V+��֞����]3��xԍ����As���%&���W����ִ�<����7e�k𫆳��Oqpp�ܽk;�3me����^��g��f5JGSP�:����!q���s��E���{���bk�+P����� |�AdeJjj�!1O�p@O(ɍ�YLW����<��P����[wm��{b7;q�����$�g�BO���D{�	ʷ|�eĳ��*Z�ݸb���g	P�,�*��@�fAC��`��T���1,�+��K,'��/ded"����Ѡ�g�t1�&��\�<�$$n��2,�냞��$ 8g����8��"ԁhCtl�����W![�۽o�i��XO���SHY�����E��b}0�H�%����J�CG���=ҵ���z��꓅ֳb�	����S�,J9x�����]�̥�?���@�=/���qZ�9ԕ޸�?
��=��{����J䲧���c�rƻI��7S m+v�=0�Ų�22~yo]�}��ڃ�㔅�C\+�n{��A6��qsM�y�ߡ��>^Z]gcڙ���@��'�s~a���g#�AD�:zg�.�����d9��	O�t��;l�ҳ��D}l���8�\ܹ�Gbb���7v%����w�+6{�����`��o�8D�\c��C�z�mԳh6�3�{��U�;5�.8��p?�<���b�2MO�v������/�V���	aAG��_Z%����<(ILN���tu}�ϼ� �զǳW2���{j�ZQ]h�"�/��߅��C[z��懑�~ɸ�G��@�%��-8�]D��̷w������~����!n�6��l�ʠ�����^�M"��҄�����z�i� �4".N�ؘ	��W/��@ژǪ�"ʚ���i;�~����?��vn������I��f�~_�~���k]�I� >�~r���zohP�渝�:��@��+

䰙�_����C����O�^�w�������#�T44� nm�"2L_��˙���Ĺ��
�Ǚ����͈Żmd���4.Sla:�T~����֪u��mX#	"L�KK��0ME�����.-���s�@��5��̌�l��t@�̂���7333Gk[��Ch���3(d,#�6�̹f�k	���¹m]j�F^5�U�>R�o
� �>}�����Ľ=�z�.j*��?e��^{:�N0��	^�����*�ľ��&�z�{�՗L�,���۩���>y�l�o诟>�������?N���`�pߟqߵ�f��|����L��"��CZ�2���t��|5_�������Ӿ]���6���w�Bb�2���?ɒ��y7&+�3p��VOv����5���$�� %�M����W����zrW@K"�y\���3�ԅ�,�1�=M���*Ӭr^��>��y՚]Y\�������)) 	�Y����K�wrb|�1ܛ�c�����!/''7}���DT4�F��H���{�(xj��ɦښI	���ڗ��,wc�&�̧c^@{b ���`s�Q�ӝ^�0	jn�I�����@��#r;�x���-���#���*::ؒ+.w�ɫ�����O"N+#}��^��uX�}�͑���]]]4n#� z㕶����**0�J~����ƌ���
g�hj^��6���G�>���q0e�rJl�S���Р܉���!E��+$!���� ܵ�������@�Y�����\5���0�Rw�~�U��e8^������=A��x^Sc.Ŕ�$�$=۪V&`�;=�P&�^����܋է���,j�����A��2^�Qo�KZX��V��v��=���.��w��������pqq��G޿���y��ɯ���O�O�d
�����a��Ƿ��r

-������xo�\X�w*�WtX�J��& �A����K�v�����!;�祓sT��.MMM�!�#�@N�8��&g:�BEE�IO:?\%&"�cqlgx|�Ԗ՞������Gw/��rNLae�e���5Ԣ¡z6��@M�m�C��	�Rбq�`[�kǀ-����B蹸¹���_����IL��t��w�"v	�]E6Q`ۉ2���bT+8��I���pH��%''��N�U~����?.�k�CI�B�k�>��)�K2R��o߆�:���d'����7���WL$�7������Bv���lzigqs����5ަ�.\qy(�ʕX���N�����'e�$�����+Y&�j��:;<G�wtdV���Ƴh�PC�,5��,�G����k( ���q� h��¹9=�9v�xV��ufrF3*���b=3.�YGKK�ήx�/d�ڑ�b�k2|5-��X D������D11�:#%�S�`�Z�ܑH�O���r����E�������tMnd����-�$%6�7--�R�N]���F��-{�S<N�h4��R�5)0ۡ��:���&�O��A:5}BC	Eݎ>+���1��M�[���S���
�~uu԰��V�5y0��㩶z��z���)�W��4mj.��w��feO��ס���B�6�����+���O���XЃ!�u`p�VV��; U���Y�Cc��v�E�Ĭ�Y�����!P������b�x� ��.���_�z�	$%�\26�_�����Q��w�.���4���^b�@O�����.�F�L�7��k�95P\�߼}˵Y���Y����_�3=�$�wzj]��Ԡ#�hc([I�yn^�R�������R��SMPTթSy;P���Mn��ԉ�ŏ_1��4I������@��蚒]-�8����e#�����<̾s��DsıoG ��¹lr�۷o��M2���""�����	��O���#:���Ui�X����UTC�ￄ���+m�� �t�L���/")i�"�8H��=I?|*-���{n��&&����/d.�>�ࣂȫ��*..����e$�� V�u����#ҵ׺hL�>c~�:���3-�_��	=���nnn���v�ﮣC{�����1bbK�ʼ�M��߿��A��i�'G3����Ŗ��D�I�;ZM���l�!}Ϣ�S85��r,��RC]��;��qq�AɸEZZ�%_�«������r���Tvvv".����/O��	Mdkd�
&@�V�i�dP�.�L�K��6>w�m��B7B�2'�<�A@������|*������gc�M]]~`��%b@~q[���-�)�^��z���
���qӀ102�(��(J9��5N�׳����P�a��x��f����(�P<�lV��v?9$Z�ޅ�r��L�����ULnC�W�lz%�K�ǳ>�Ꭶ/|&�/^w�@p�4W�NU0D�iǡ�{ ��@@�Ji�����/ �BAA�t�>N�)�am�AP/-e|RRhR�n	Îl�UE������j@"��(x�z�v�D��tvp�i��1a}�u�8���qEw�ڗhX\��"�'@S���|3���;�����&�Hm�0Y������b�|b�m�L�����0�~��S٧�;	��v&����+l�a���W�V�[*�C$���S���S�P~��~��粧������1$��_Y:���?���ά[>�,��C�,$$��	Ǡf;y�0�'v���i�ť�H���_���^J98�T��=i:�1 f陮H�qɼ6���U�`����������ql0��%�~4��I�b�w����Г�y�����Q3+��A+����"!!�<r[�FE���8����NL�T��z��Vݽ{W����r�ׯ_s��P�����Hݡ��ө��AF|4� *�*�]z���z{�S;uh�C�	Uۀ8:��M��%aX����	4?��]+���ۢ7�K�Pl��u�x�-(�΍H�?ռ�����{O�Qx�p˾�� 3X���I�XDDD|�t�;�!p�)`�n=N����+A�&����ˀ��1��h�[���js�dV6QSJ�O�P��T��&Zi(�j�b�+�v��_d5-���^*��40����x�P�)��͡�i���4+��<�H�s�?awo\oVv�3 �y�w�.`���kor�fd&{��:�ϑE�GI��.���(O�hJL�W����P۽H�;:�Y�W&;/D(���ɵ���e���=}�&�9£fe)�~� S�I�G��7��g��h��ju��ϛES�F�@Pd�����~����X!*��Q2�$����{��![[���*���~���O(b�_�����G��k� i�������+��r5�f��<U	5Dx�G�:�aw�ʞ9�k�8?�ť��3���G���Ņ�n��m�m��|p�s������ÎeeeD�цX	(-,>�b��?�������>驄I�9�^P��ՙm�0����LP  $�k�������SG��e�q�&��X^��&�cckV�o]qq[zBM虙3SU[^ͻ��!=p��O�H�{v����ʄ6�p��RBϓ`,�YYr'rNJJ���%ffm��NZ��g*%�	���hhh�1+�~���_�q�������v���i�Gs��/�aa��˫��J���<4��C�񐃃�_�?XCz=;�F�S�%�>.6��lO��+��`��b�m�ʊ�{
��*I�NJ�������Z��ӎ7�������n�5����s�qA�BL��d�+������@�ۮ�5�[��3�Ξ� %]P9N��%a�Ąx�1V���QǏ�o}�A�Yʤ��"�rH���d/�r"��|��o�!%4j\�P\|6�`?a��_J:��g��(�����|��u��?�w�&!B��s�z�oѤ��'�5�~P��N��<R�$���Im
���t{�n�Py�j���b��a! ��|/�"�C�N��2�-�D{Ⱥ*@�W�����͎���[9Ðo�&���٣UjA;���X@,�}
?���l�m!}��Sf>�RV����ޞ{csFJ�\������zڱ9Z����m	u�1w�V@��<��I�t*��0翉nC���qi9o� 	�S1��I�<�w�|�JRE%|�
�n��ߟ�2;K��wD�22�pΈ�	EP��(�k"�p�	P�SQq�=����+ǟ��Sۇ�xb22?��/�kΧ�*::!»�ē��B�r��YY!UG���8�ޟ��'kz�81Gi]Q\�g��"b���mwU���'�`G�C�D��A�,w>=�,*���Vd�Aԃx���\�u}C�ȂC~]sM&�)	���j�c�V��Vaqͬ���٠�.נ�ż��fP۵��ƹ�ޞ��ָ����4&��4�I�c�����ִХ�qBa�r�ݎP:Y#�t��:`)=M~�St�"Z	�{���TM��G��Ĩ���x��$/�W�>Ч���KsŔn�.��D�6�j�:�����؎�x-��m���5X�~(K����0���s:��7׫�O2���FF���q��QU5�ߗ�F@�AEBJ$	i)�K���)�n����4�����z׺�@�L���=s��� 7'L��WO�<���937w��xo�ӄ�N�,]�s��$DA�U(Rp4�+%���0WK�&�޸q�j��^�
���u���CN4��$�Oê�U'^1�#���7g�� KK��Ȩ8�;<�å��p�!7:>�v�X�����M�{�&|��]޷��9?wP��"�]�����0���l�P T����%�{��1F	D&!-�G����ӛ߭��� (�Sa���e�@iu�y������� !̿q��v�?*�NZ�����#I��_/�6�׸�W�7� !�T��45S���`=�D�8(֦�0a4�����ȀjG��XVV�S�U�_����Ә�&J�i���..����{ KMΎv��-se��~pQ`���0�_��$`Sb�8$�6�s�|q~�Us�
�V;�*z�z����E�'�h����Kߩ{����}K{�f��fKB��&��������l@R�wd��_~����r ���IAo<�g2�����ii`�W����p��kR�س�>��� <z��C���=C���=R22��5X8;7��X��%l���v����D$N��r ���k��ދ��|��h��[�S�}��d	�w����ɑ�Q����g��ŧ�1t�&vN�a�r�=����9",w�{ �MV_%��ƾ��WD\�-Y�y���y�cv%;I��*qY�������@{	(0�$�zc��2ʶ/:C3���3�ÃZGo���q"6߅Y��HFM�[e5:�;≁�1\`���'�s�����3�2jO���r���G��U[[[k[[>���+zԋ��,�D�V9�Vz��,�^�~%×2P��6z' �(BLC����b%�Ұ�h�eWQ�C9�>`��$���v[�L�ܰ��JN7���[ṫ�������w�Y�o�0^	c����~+�bM�#QQڜ�.�ck�0��?~�<h����@���Q2	�Oj������z�H��B�D������'zލ��ڛ�����(�{os�z!qOd�r�ʚ777h�bM�C5��=�r}�I2�t��k���)�h<���J*bN�C��-����?���8~�D�}�ݯP�  UL���$�W�o�U���6�il�o�}�f�B��0X @���x?�L���eJ@���K� V_�ش�SV��,�U�3�(f���_^<�*�n�ѷ���k�<]"*=���XJ�(��M�&� lXf^^�,����ŵ}��~v����[��N�����y����Ui��p31�dee�Kp��a�Sp�X��kaR`�ѣJO_#t����+yW0�Mx3Ktb"A��]���R*@�w	��3A�,���ר�P�&�QYIK@@`/���{�/��u�~aCӃ��$*ݾ�(g&�K��O7�x0���<5���?�2���e8�E�{��H�6=��1Q�ٳ��bԗ�ǋ4\���H��_��(n#*�($w6"�O���-u&���WS�jem]ߓ��xAK��uy����5 +����C�Z��II��J��{,ym��V�_"q䱏��p����^!�*�ʢ%�"]���u����ijɒ@��u&�O�'Wy�@ ��q� ��X��z�dRW�%�ܬ �NV0�e!8��LF� ����f�u�7�1���Afgg�[)TLm=k�BN��*�U��,��+r�����ư��yFV{p��E��M�����Jj�����6tpd��&�|�3�u�wA�����s�SP�%w
�(~O#�H��NP�����ʃ�>M
W���/t^������ ���/��a�������N[K���Dх� \��)wp�H�w�o�ՅM�b�f�������� ϼ����߿�t���7,v���I�����i��W��� �CF����>j0 ~�7Iplg��	�_�
pw{ip� ����3!�O*�s�
�QcT3d�����Z��ŧ�
		������NI��d!Jy���&z��T���w���V�����\�%PI�6"��ܧ�*R*��<.n��d��D�K ��K�Eb�x�� hR���i�����\؝��e�m�&{UnY�^����
nn��q���R�C4���d�ɋ��hg��x1^���'f�<����X~Jt����U�l^8�]���F_ϭY4�M��A��7�����{�,�>QW�Y�M�Cꀵ���E��ԋ���̼��.w�����"�B��O��F�Lq��Q�B!��aa2a��4ef.�{n�O�.59^7�R�7Q>L+�WA ��������o�7�[b5h�ٔ��v�7A{,|�� ��C�I���ɃF�Cuu��U-�xP��'����Od��!��'6±�/|�6Y�/p��Óp]�m�w�xm���AsAsU�3��c!P��޽kH~%U��1ќ��S��͗r��դ΋�W����("��H��r��Z��x�U��v�H%�`)�����>|_I';]��]�ء3Q�rm(iq�]r�2���i������vS�t�k�@��x�)Rh󽳹�%��,-37�|O@�����zka���κ�TZ䜞Q3�I�r�xzzz�Χ��w�7x����p�i��r�l��|i�Ke�Z}�&�S7�h)E�P����O��[�Ptw�]Վ���6�p8����]���~NG �MQQ2��\.󔆆F0��V	vvL��u��΁Ǚ c�}v�8��y�홸glX�}���l�4����&xwE��8*.��>�u,3㨫�+=|����r�YA���aj�A� ��d�Y���<�u�@��M����}W��X�j+�{�����sg�O���m&_���7.�5�Ӻs떌��T��`�{���s��MIޠݡ!v�f�&�-�ˆ�`�� ��m�a��֍�.z'�OG�0#����iY"��1�W2��L��Kvv9��h�F�m>�=5����SE~�`*@��=K��揢"��|S�r�Rt��p2���􍛇�}��ΪWp�,C[ɸ�
��L��k��N�G���*775�۷o���o�8�'O�D�^�y�9�֢O���C�ۈH��1�������Z�џ?ߊwM���V�<�
�qnv^5��Q���҇�Sss;Y��;:�r1�1�n� \�h���'�'�6�YZY��"�BcbHyB�
N��?~�x��	�X���p/�n��%��j�U��~S��)57tTn����Y�H��$�pK�N��~qcSS[���N̺zz7�Z�+��\���@IƸpQ��$���������,�T�ax���+Q):jR�0!�� �J=�鯘=�ݗ/@��� �`�C��:U#�]5�XFu����~�N��6l��MX�a��[���@��e����ۈ�h���#�,���]֖��t��a���FN��[^G3�;mɭ�@MC�eǺ����ΪQ�f�T��
���0Wr�Pk��H{^��瘝ʼ���H�&�/����%��uX��>$j<yo�=,h��0)ޒ�����=��L����F"����o6���8�j*���\A{�:9�x��rr)��� �p�B�Mn�����m��e�9W�n�%t*�0W0d�J��2[Ԁx;���k�4��@�t��y�)y8�㴴��{������%�9�5#ƅ#�^�8iG��F�*z�moӞ4��>qW"��-��Qn�N=t�P@P�U���nG�����n��ט%�n��L\����kpXsY�#1�oO	�Ys��7dG�-�oC�~qNg=���ʪ�X�Т�)/�;6�bgb�۷�m"i��RR����g˲	➽/�*QG6B����;I��Y��N���N�_�$.�!�Pq��C�Ž������� ^t�Yp�gQ8L/)*���m�ρ*��ˈ�Of+���/��g����G{�ө�X�=@��[�0c���j�;az�����w[�0�5Z�顀D�	����
�nD�}�=��b��h�����E�E��������j0����E*O��@Lس: �f9�򃟭�J\��e����ļ0�p=<,�͔�?�_�$%��� }�P`����{��|�	r�%���<�*�����'�vvw%�vM���K�-��V�qf4��I�Ύ梨���mY];���*�g�}j1RQ���,<<D>19�12uqXR��CG��dMf������(h�9Ď8,�J�X7�G+���/&=��]��aZߊ�gmm��s�L-Q0&A��C�]1����#�bQ830d�d�_a��(�  U�N�A��������=��W�}HH���9���j�ƺ�UJ%��w����@'�$��쇶��'Ч%A[���<�̄h�(0sss*�)G����5o߹#�������ɰb���T������P�!�H�S={�t9-|��oJj갮O��:�5��'��|<8�2��kW�!<e�2YHIIͶ�K����3��.�,f�$eut��i�� M�Y�Z�3��%�4��p}7H& ��H���s�h�b���f2;�<��.|�6"BƮ"���p$jt4�� ׈HGGtVkM���\���d�1j@���@@��/�T>�0e��hҐ>�$Q�/N�!�^�TWӳ�_	����|����o�ȿ��U���"�[�wE2��n��h��L|f�D�lVΩZ�ؽ?2��[�@��w�آL�.�U��ʢl`��;0:�
�4��D�N��U�u����/�L'���0�k�����8�%7�.ȉ��<�-�Η* f� %6��\Ej��_�x�+Eƫ��_�U�>F���pvq!���+�H.��4��ڣ�+��h���W�eH�KI�z�c�ט�|�S����}���֋m��D�)cGV��(�_�K�E������X6rpPK��ዩ6��b,��Jw�G�ba���7����-Q�V��.�fVF�y��$Ǳ�S���{��P^.
���������ˮ�HB�K"i�XJ|i�n�7X��ZƫbU�� \v[R�^!]ݹ�����tl
�\M�~�2d)̗>|���������L܄7���L�bӠ�X�MYY�}������	�l0#v�*�Mp�1��g��w�<|�]�	m2�2m�;�]� t�G0�%�	C�����f�j����s���I��������M,"z�g�>@����ٓ����O�i�����~��FGG�;�
��N�#�q�{Yı۾�G^o�g�ϛ�ڶ���T%�z���o����d�������ӧ���VW�w�F�U��Q}kBŇwz Zш1`��hl�5b�_��� Q~\࢕� � q�F%�s_�t�������o���?z�h���@�0��*�ti�}�U7��.333�����{ T���u������'�w��~�"���I4��.��)�r^������JBC1���x��Y����\o�恅�uQ�	�M�uq��G�S�� G� � ��Fх�8@���Bn��q��m]bJ�] ��wމv��x������������%�����O�.�f�y��Wv=�������W]!�י��Ѩb�n�>@a�#�φ��p ��~Lt㪱����t��xk;�4v�WzK+��]�q�!�}�Yt��:= ��\�탆<�\IP�~���,v�8_K�~�����<�k�G�&�&�c�����ѫO�>��I��	��?8}��B��D��/���n3p- ?��(X[�XO�4}�G��!�V!}>!�:��� �oQ�� o�� ��cN�Fq���R,�i� �x=���4�gϞ)E���̴0��ii}��M9v6��]"CTQQ�jN��Z��1.+;�hE�tm�/hZc�����j��ȗ��v��~K/A���Y�y�~����7m��)Ⲩ�1��`gפ��??<�Uk�H�݅�DOH�5J&�h����&�U/o��h����1*u���Mz��msB��8�u;w���*�*���w#iEz{�f�a$�=�A�R(	�;��K���Ŧ��iTz��޳Cu�!qy���� A�b��(��[���풑o"��b�@�\��mY�i:��pc,�eIաY�������q��X>��o��kiQXt&��HMM�:gV#��I���&�O��G�F���^u	Q)C���:�|�y
w�ԫ��Ք!u��]p��kn���.T�G�C��Ru1)��=��'kѱ�KWM��?x���G52T�J������V�����|)g''��*`gm�������V�_��Ȕ�`�ta�t��D�/81�� �(�W��ʑc�B⻭,��J�*��h<���u�"��7��I�E�}fc?89$�A�"ݧ����)����ѣ�+z� �di�@���vyq�3j��֙���܏Eǡ��8Zl#&���Q�!0$<F ��Cޗ��<Xו��}L����g�{���B�wՠw�x=��GD���~����N��s��,�tW�����\5��EOOO�KsMhA�=ІT�q]F����-r
��J���G��b�2ԲD�"1܃�g�.�������|��#��	��p�LKCeQ�\ﯚ�cgbBqY���idd�;����s��F��k���~G��_,���y�x��ۣ�F	��'G�	hx�m��ɾƯ;ڙ3_�N	�
U����@W�	s4�E�wzP��:kB�K��k�����s~r��aaafp���� 2��[��
F_�㝎b�Sec\�:�Ǐ�^��t
�����h�)�,���~h��]`:���Q�o
��2t�F���B���%�A�{K��=J�Y99�G(�ξW�tZ�Ɵ��c�����P�\���	~�6X��c5��fff�ՊU��P��ӟ�����ثc����GfN��2�N�����5`��U|��6@̻@g�����]BEw`��9?E��
V��nv���YFn��״$9�I]���+�rpU���\+4�G��
JJ�y2�Ń��{@�AW;d>�Zn߀���v��3mm�+"��¶��0c�*$�B��<����aĆv��Ց@aA�
@Ã^VyK-��yܢ0��r�[1X�|�Җ\�9�-�_?JÇ���Sr�����F��]���v�D� &�v����O�0 ��V���5�gZZ���9Zs�_�渗k�#i�'��n��h��v�+=*SC��&ҭ%�&r-�Xn��P3���c*~���v�B��xD��o���a?�m=�M�EVGR�P$�0��48(\�2�41z�愰��+�IY�J���}��*�w�oU�U������2XJ��ލ��#\�̪|�6���!�K�K��Ĵܓ�����O_���d�4��E92��♦fY����$zZr�`��w�H�p��6�`E7���el`�:�p�-�G M�=v�8Xz����Gi=�P�/è��Ĥ�~����w���_�P������7["�4�$�?�`cg�LW��D�`e%cg��l"�d��G::�MFߕ���K��ϑ=��Aj�����I9 �\,:��@^�<��J	PG�A�ehSW�aigW,��k�
��'��]8&u]й���f�;||$ }\��ji���T�ګ���˃�֕m4��L�! ݢ�u�uW��!s�IBM��:��%�x=�+++W:�C5�X~*N�g�.,,p�	�����@�a/�L��%�P�Fi�s��V]?J�V��%`�d���!���]�>d O���Լ�E�l�(�Km�wl�����9��c�1�1S�<_�o�t���˼�+�}À02���BzBFK<qD ^�����h9�	�ǅ*� ��SRj��-�w>��,F@@��
��	U�h�\���]�r���NUW��6&�T^s8���'l���ҟnzr�*+jV��N��}U��7���'_��ls���j;$���K�0���".%�iv��Ed��_!	���G���,[rc,�<N��K����[&���&N@>7�a��ʝIQ�#���Цן#����ȯ�"����y�[�񰉈Zң9�
	����,H>?{cZ(0VA�{d����C
�Yh�󿌕�`�uN�X�M��}��K����E`m���o6.\|J1~�m��N�}p��$��Q�f-Э�!�;<ϟ?�u͜�ps+��X*����e0;,�]�0�����ǔ�*EXʆ}��ڠ'?��H�a� k�����Th�qK�=�$#W_�Т��i��Y�Z��V2L�������_7�}�U���b���A�5[��˂��2��Â��%���]�.��H��jV���p�������L`�1��v#��R��'U������e?�{y����1P�Ơ��:*<w]8�.�m��#�<���<kA�����\-����N��/�uE�r�$�364ƿ�G��/�C�bb�o�ٖ|���{F.!�b*	��y�g�|��o� p3�e6�Pv#�����Lc�:T���7�/���>x4��,�Q����\���u��˰���%ӭ�*::�|�V_IiXI�F�'��W-���b�����f4y�/���"낱�#�55�L�K+'3ʒE��Q�W�qw���=Rk��ȡۯ,�g� ]FZ_?a�h�:&z�r��pbL��	>~�ȝWl�����+�ڈ�s�l��[",�qN.�>s];�M	OC yq�*��vAa!��',
�j�-`� �Q}�dॺ9 #��/�bѮ�
����������O%L���mgppPub��z඀�p����C�)�H�۳��Z�����d;Z�����5�����|�Oqy�(t��������-B�1��_@����Hx������k"nC=�p��C{w�|���;������y7>>
���l�Yh�M���Y f��>��{||<Ծb(g�G�#Ցl��4�����K�k6��D^��&|m}��yyy�����?�\0aW�R��x�r��!O{{{>P\��@?�B:	��|&+=�`̽���/�����u�́���ϟ�LK�l�q)(�W�?����_�T���S����.\�9)h�ި��ڹ��;�t0/�ɳ�8'��"�1a��%�JZ«��557? Fos�|��3�Umm�44޷����v.�a֦�c�܅f�������5o��wn�%;�f�\��oR? `jɒc%@�Q�1���MFk�%��S�J�A��6㼟?�)d;���EB�(�hڼ?�;�<�>fk�
y7��5k�:��HN�{����z%YU��Q�ԣ�[!H�T��N�������%����wR�̚-��z��O��!޼��ִK�M_,�N��o�\�q5�"?���&�'ߦXR�9��O*�WO]�0z��d��/�����p�#n��aܼ��?5���Ve��]�L��<��ۈ��t/��_�� @l�h�d>SL9�g�̗|�,�u�v:)�O/N��D��TCG1�ա��.G$�痂%��w�VX 45>���seyy���m�'\�'�XK2��)b�I�i�׃pt�8y{���ms�[)C矅M��mG�����|���JI��M��K�3�k)���D~�$T�w�{�����v�6��%wW�R:�43��xX��h�h�a:�M^<��B�wvn�����,�����#&Nw����ѳ�xmP�z�uڰu�űl��T�{z�ZZ:�O�����P��~���D�d�8��qEU�+�+��S\�伥�tJB���6�(/����z΂ǹ�>����9�)��n� �Ûc��R�b��`[��Bo�����	��99���i�V6���OV�A0�py��ƧN����ʮ.�������b(QY|E��l�i﹵����S�����6�2���Z4"^�� �T��^��e��{�@*Ԇ{��Ӡ|����ޫc=�������0���_~\�y)`]XDGG� ����P>�ڮ��Zd�b[�I����'�Z߄�)v%I�/�l�a��'����$ �����~G3�{[rH���l�$Ď�U������]�� ] �3��i2^�8JB�	ҭt)ɛ����Z���e���B�X=��z8'���R��כ6�?�ݻ��c�ڢ���3��u�*ڟJ�>a>�3,��gϜ�ȲP�Ҋ���:1 �$�<D����{%s��v�9 7\��tb�����K�f�Mn�q�~~��Y�=L�$p����˷`~�?�����5c)��6-���8��?���ԏ��l<���������X)��hk̠�X�M��'�ڙ���?��R	�C����
��8����g��aQ?X��X�H�SIJ���v�O��*����oZ��11�bKeKI�NN�`9�KK�_��4��H�&������U`h4g�\:u���*`���n�mE�M��/yb`���������<�P[.��~.C�ũ��NV>�i!�f��� i�5��О�4����k'<�������r���5�1�mf��#��d��,�@R����E]��]7�*z���QMXޕ�
T����|kt������U�ɉ�f(.���=�*i��K�o����y���))>f��Q�l(To�����E�R�/�sPFQ�ZX|�mYh�Რ��&��zϿ���b:� ����V*�G����}�f�Ο?�i˽��Bv\\\C�Yo���8X��[�x}ݍeZ��C3��W�f,Wm���cJ�!((ȝ�7>��n췛+6]|���,�s\�����<��k����r�0��f��,�� 8*6+�T[Z�#᫪�..��0�5g����M��sJ�����X9�begt�u�����(��2S�H�܍?������Iq�a(�1�)�Ӝ��k��f��z��H��£+��3l%�.�j��8S�H�Д��ˏX�k0����\�F�^s�u15���{Q�g̖���5'7���D�"��9>Ԟs�Dr��0�,��©�om*�^�ȯ^�~�5Z��ˣ��<�V8�S��{.��OZCC�%��&�"9����]���bלC�����H)��/.\���͚K�u⇑�ŸS��TӑPAJ^���w��c�%�[���|��)F��%�� �	�˭،����}�a�b���<�s��|����E��Ye���[X�`9�G4G��gO��W�C���D�3�X�T�����i���s�s">%�N����� ��ʊ�z�\�jb}�U����Ǐ?���ee��7Fz�ܷ���*�ިTf���Y4�� I���9�'C��3*u����z��nƺr{���ld�#��aÌG~�����O̝c������;ڼ��&�@� ���3��X�B �[����ͦ��)b��[c%�)ʉC�"�X�����_�ʁ᫩�bP��l��
�����TMMz:MT\;�m~��]r����F���@$�c��/�����U�%,KP�w�����ڂ�����kۆ���͛+����S���%a1�_�8�[��,Q�8�oM�O��{�͢�ڟe�=�_O��-�Ȗ~�m�ɫ����Ύ)�Zi�� �|ϊ([k{�ڲc��D��+���ï��@�-e
Rd�<�Z&��W�^3�S������wF��{A���Q��vv��X�=;���pn��_]]�ׅ.��#@	FQ�DYf�ȠDw$��6;����s]˔��۪�{ٵ�R����M��������?���c�B�\:vZ�?�tr�t���Z�=^�����y�'Рn2��>|x��������_F�GGB��NNN�������l�,,���v�Bo�%F'ߢ8�l$��-G�O�N��t�./�%��=b�@9Z+;D5/4���=� {@�M#�D�c��h���(\#�B㎮��k��3���$$�X��(���-�쪦��0����ҁ��U\�p�QR%Y�<h�����nN���4pP9Yiю
��K2�.'J����Í1��p�A�����ةq$���1��m2^�^_�1�4�b/0�q,%�>�N�[{�[�U�6���B�{<����7�T63㨨�O~Dpf�1�r�X7�������W0bE�1��5��Q*pX��䀌�8�sF]x@��ϟ@<�=��ba �Mb��uv�@�Z{�.�_hh^,�x237!�����߾-���"�������~�z�- ���u� h��~�1	�S��zO����3����H&�Q��{H��<�Ú�-U;����i[�����{"X�ĺ��8*�o�ry�"J]�|�X�X�Sv�O�%v}�����$��Y��-��@AP�7�P/%�RNϬ���|�o���<'KDo�xM�H�.sz��1A����F+(M�Ȉ��M�]qt	�{z���y�`��|[S4�s,��׸8�W�^)E.-.�N�NӃ ���P^]���>Akk��s�����5���I�w�+�@���-�����Ո\F1���������RN߄���ޘ��{��eb ��SNX����p�z�k�˓�����PB�X�T�x�e{�D�{��X���c�� У+��s�"aJM�	�I<��c�ǎy��޻��&�DD�,���'��y�iK$th�9��֢/����l'�-h�5��S�3�������2
���'Y�7�B��ژ�;�[��yyi�����z\�� �eԘ��=j�w�*�ᦤO�X�8�	����@�$)wc��\:<�d��@�$MK�5��c/V��D�;d�&��ƞ��N��k�1-v!'�8oK�;S���8 ���O �dk�����<��t3�s�t�fk�XI_�A��
{i��ـ��O��ߴXD�(V>WE�E!�{�\��u�(�_��BL(�9�c�@RF|����W8��j���'�#�,9v���o�v��\�R(���p}�� dPR��
q���u�Fvv�l��媅uE�S~k���~��lU����eK*| �D\S23� )��n�@�/��)��N��{�˔�`��{ M������Ċ��Dt�M4����.t�33J+�&��In��m�ɑ�˼�����q�Q�4��������d .6[L����1�A���[�Y	d3T�J����`�S/�Z*�h<N�`��6�����8K�U99Jb22���o�?�L+*z�a���5f\�E���p~z:�4�Z���s�������Rut��H}/2���1�����J���1y+�:���t�`s��[n_Ns'*h��`'�4����z�@��ٮ�Ӟh�����wi�i�?u
�� ���~�$#ADD��f���\N�����XA��� � h�~V�4�gp�K�P�A_���7a�U�K�=o~>X�B��r�=�68�$����*������ Q�u�(K�Fߤ����H��P��޺3$-���;���Vf"QB/>BYEZI'�DV�ՀuH�YЈ������츻vF�i؈�k�G��#��=�����<���X@�~�x����b��D��y� |����ݪ��F9r
�?Z�Dr��n-�O�ZZ�,͇�M���a&F=�Q��Ӓ=M�`��9m3cВ8�8j��5�֙E�Nw���O�EEE)߲n޽�aie8:l�~r��eֳۖE���#�������n�]��U:I���b�3O�i�9�K"LI��������O�>u����P3�����򫬏�Զ�`�3�E1R߱���A��j�%�t	�Zi��W�q$�+���i�@q y\l�]�[A����1A�=��$�P��'�� ��� g*�FMM�����E�i��-o����Ѱׯ_�u���b�	�[
0�<O~�Nb-uv���R�NS�vW����\5��$=���W�h��ZA�>Nt�ʲ��j�A��DL��>u��qW�R�s��p���J�q��-������H�]�Y,(�����]s�1;��G��ܟ�cب��I"���ޔ�_죆�2�f�������#GW�����)�h%?��a��b Ƥ�9��h6)h�J���0''(��U?:�lMV�o�O2�bb{|��)}��ZZ?9}`��
���쨰]wNn���)?�H@���d�)ݛ+�9�,m-����y��b9f�{�b˕fjJLJ�����տz�5�x�;z
9�߹-)����^��S�{�pӫJѝ�U>�������������%��2(M��E����'E�ǽ�n�����Bo�Z���wb�V��I�LO�Y�=ݺI�������:�2��e��pk��*8x����w{S	)�е������ņٚ����1���lL[���䐩��uv匾r�__��8�ki`�/�8��.�<�A�> �[��ds�p��_S���#+��Fԕ����*���7RR��~��㆒��"Y_�_�$�R�Ô�����b-��<Oj���$ N?�{Tl3���\��i���A�2}�R���s���W�Ga����۸S.�M϶u��z{I����ت��M�Gb����;�0�1���!Zf3?�����;�p���Z��'�W�/�	�Yz�l��>��a����7~a��RA�@�PQ��Φ-ʶ��׌h��|��{w���?��P��nP�g#eX����aق:1���׳�NH{��J��JS��}.yu�&�al���{�d2��Ď�8E2��
�ք�e��4-��F��{���,�H��#�'�A��y��b��5}��gl{y��3�&h�F��Whh��Oc{��)������ӷa��5=eq���<9�0)BA���VXP�~x>��1a}U�M5N��L.�Ւ�qK�]o2��H��Z���I��0ݵ����mpڸ6}|��.c̨�ݍE�� ��{��܂l?v4d�_�����Ř��>A�EIs�؂�M<���H�o���"ai�BRQ�g��<'XX|��c[�V������]].�b$n��]����?-��z"'�|���@a�1s�E�FN�c܆m3~`��H�l���:8<�j?�z��|Ú
Oa��V����j�fI����Tu���\�-�l�H��ڨ�^2�r���:||"�O�U�����(�ai�w����h�yyO�>��$���}I�dvFY����\���b9�~⊆��*�����g���h��ι,��D��\HT��l\\r:�S>گ�������ni�X@���s����\*���靈"���7��2�����^���eo��+S�Ħ(�lda����1�#yh�!����[o�������E��ڒկ�t~�=��{n؜_�#��OBd��$`b�q{�=h�K��\�������������9�}���*�V8'{0/��UP���%'9Rɦ{�
W�Z��Eu�l挵���kI&�{#�f�j����|b[-�Jw��>�~��R��<���D_���17u2X�R������%}vIE����T�k���)yR8 �K�ִȘK�h��h,,�H$J��}�"��h��P.Kl��"�oOq��[��2��T7��*�\��G1���n�/�>���m�|�q��x��)2k��Ny�S�X���+0����|����ʝ]���?�V)��^}^�J���7��Z�G�����<��x?�S���|�f�H2]"�cv��;��R!�{栘a��{��)4֧�I����{/��������������p�7:��{c��o�n�H���1��@�4����;Z�x	�.(.Jd@s�Q���`4nB+O�l�v
֥Ʃ�g�<�:�����מ	S�i��\_8KY��jY�ψ
�P�~]������ ��TL�4z�i��CCX��=ϲ�έ[���ӂa����g�İ�=K��c��d2���ؘ�C�.n0�����^���p������P�,`���?
�ք0ܷ���2���}fk=�����|o��L��y�m3I��?r���b�n�K_mY����Nz��̣r1� A���lV/�d�KV9�D53��q[����1s&���>��[��N"i-�$��@ȭnm�v!�/���r����Gi�����jˍb���y�-%�*׸��E���r��v�^�ME{1�."�5�¹���Ɠ�,ySQ3U���F�� ~��qd$ǵ���&r�k&��P}D��P�(��&��Ӛ��`������MVk�qEF���z����)��Y��_���};��Q�����ٽcΏ5"s��8�K�-��09̎�)�F?�	�u\:qafF�ʨ!�A˛r�sL�-�5s���z�����?�6'�#��R�q}qV�m	~��QUήun'%[�[���|Y1.>�'���M�1� �	�I<c��);V����u�bp��$$n��?�	�c�t}����i��/.�˽�~�Y<�R�Mq��_��\˴J��b�c�����>�-�9�#�k���J���6�0��{���뙔��Ta�@j������)�P��l�Oo)=�iiuVs�~���qG���M�t�"�=���{�Q�@��$��ΘؾDo�H����د��VO�o컊Fdu4�7!��f�嬁?ǜ��w�ݢ/=Y��8�F��'���g�t^�c�~�W�<��+������/-�y�'y �D�~��	�>���"s�
а����D����=��s�bt��(�U�n�q���@ɐ���e�+��n���S�c.����w�M���w2|�_�v �K�}��g�C 1���k[ݲ����+u^y���'Z؅�rw:��I�3��W�-Ό
2u�w�7�����:�wfB��e؉�0�<,2�ijw����.zG��LH�$^�A ́��-�dN�Ӭ�Έx H������^ָCRU�G��!�=�J�,�^o��yyD1� �+jN���z0������Vګ:�x�I��177����������OY^��|����75^)1�eO��]6�R�S3����R>�rE��XD+n�*GP]��rқ�5)��������홺`,��ϻ�����"���R�GT8��.�~����C�E�|�L�0����e�q�5BC㾒E/�ؕ}�q�z'�!�C��tb��ܚ��ȿ�1��č��b��(xG!/��a���ڧU��?�[��: ٕ��u���lƟ�l�A����|$�w��/O��Ξ�q��Y�9��],�r�+^��a�z���Y���ڒݚ��h�d�]_R�S��@��	%BA{ق���iY�r���^��N��h����t,����Om��.�䞧p>rc� ���,0�Dv�1�^mzrc��D�����(��N���K�CB|*ɱ@�%���״��`�e��ڣo1 ��eo/#����cB�����#��������*耠b��o絺�N�2B�|�+9�~\`�	(.Kl�#991և�^n������ �e@�����wS.�'Bx����<����d�v��.�uQ�v��xU�|�h��8��A�@�ݥY<A0x�K�+sA&�Ɖ�C��?�*�Ԧ��)[_ês#e�>(�s9s0���\m��c/�1� �+v�h�܏qocv<�%FKEE�hg.`��x���vX9�{�>��0��5���~$پ$l�/��U�@c�		�ftm��*7��x�*Ĩҽ�ڈ�����������y� % ��*%KJ��t,H#��ݍ4�����Ңt
K������,�!%�﬿���'��ى��cΜs��AûY�=���YB�N�5�Z�EbaÇ� M7C.�����#���mK雸]u�@zw��V~9�� ��o�/{gO�"�zW����^Z����7�_�K;�1n�f�f��D��]R3��@��9��ݻ/��6]��*�ni �޽u�k0�1/�${�w��8�t���> X��#�J��i ��,�텨Պ@֏�SqK4�r��jP@�l��O�|���#x��Q���Q���-���ɖ~���}�K����qi��B]V�l�a'�oΘ�3����BW���]�Y�"��
n9s��}��ܟ��B\CV��B/>#�?�޲jdϷ��
��w� �G'1�ð�up�y���ڸ����c�R��YB��W]b`pi���D�&Z]m�[��ꐼ��9Ց�
��ҁ�ӯ� K�o�C�œT�1sC�p��u�ط �byyű�H�w^3׽mv�_���gN�(��P�
m��/
�
����2,��H:�4Y-R虨q�b��6ה������B ʘ�'�����ː)4����. 0���� -;�������F
%� ��z��zM��H�����u� �iǓy]EE�.i�y̫��Ю/K�߭��(z�5}�/����L
:��\F(��q��c�G�Y'I���d
�ʾ)J*�ꖖ�����1���l��9��q����݂i ���-�D�����B���/�6�N��`�!����ct��55��g��|��e�%�Fv�����<��?!�ۂ�
7çX�̤_�H�EcĄ]��R�����a����g]DV^m���UjM�>ҟ�+���	��h��l��^������n�M�]L�+��lr��3�1�TCh��b��v�-ʟ�`%���U�������>2-�%��I�m�c6qg�̞�L�^f{���C}R:��˻5�k8�-�(��:��/�8�<j�a 93tN�V��;Qt�yrر�E�W���`S������O�շ&49�þ��޾�" ���8���i�n[��c�E
��u�K./yT̀?
["��C���Fv ||�'��xQ��~ݝ^y&%
�t��ƞ;�<�^2���ޭ;5j�'���v�VW���gY�}n�PF��vod$>�+�޽����� -3� �h��LŇ��G�	d�*d�;л�vz���ptB{ƞ��ux�H�\Kb��B�;�}鬣���#�	���oK���p�eכc�<�Hѱ<��De��7�aQ�^�lU���D�U*�/#�l�ߠn;�s��?������C 	���da��_#4�"7?���G��v��VXw�+�s��=&�s|��4ٻm5�y��=z���u���������K�7�+Ӧ�?$�Rw�X#Xi($!���p2��G� ��]Ad���&��s�2sXut� ��L��_�K�Uq���܇5�{�|�����V�M!g������Ғ(���(8�<�\��blU��Z2�@�'�x�b�篳��������n���0+)4�\�`1n�3뛛�į5n5�^MS6	8�4��J�<��K2�B��g��j�0=^�V%W�̔����H�DBO���޿����^prz�&�oR�91|k5���yUg墤���4H]F���D+D1�aA��]��{	�_��)V�!�0��3�[vT��"Q'08�@&���4Ĭ�`�ƫ�6(wr;�6r�ӄ{zf���uѡ�Ɠ%��$*;E�Z�jC�� V��\�Z��r�<\������[)/���Z��ʳB	��+��OHm�t5౭=��3��7������LgnÛ������觰-�8)�FCJ�����(u�ھ�����8�:sscX6�I�re�`:ܪ �^�&~��J��.֢Q�\�t'�d�4_&/S��u�%�/��7�~���4��K����H<3W�jO��\�(�:ױ�Ʒ�$�������d�.uQ?#w`��y�n�C�3%R�W�6�t"��}\# ݑ�w�n�gkH��>�f�P�$��j���%�|�(Ҭ�,����ܡ�i�H�4X6�omc�0Xgs=��e
M�N����dR���+$��Ҳ�f^hG� ��|ʞNN9H�ܵp�4y���y5
~=ɣ�?</p�`Z'P�<z�(���if���(h�w��H�#��1�a�U"m�p2�������g>��m�'"{�8YhƦ��ct�$;���������+��'�T�Ro�+*͟k��Z��Q�21���_Q�r�\,x4��d�>�������eV�!f�#�rq�Ə^����<�WpmT�,;KeNnLfr'��j��6���}��oL���U>��O��!�l�e��?��ޏ�d#G_ѷ:A2�7�uTh������K�w�Q{0R_qYߣ��Rc���������7`'��goF���&ߥ���a��]Z��,���>,�N\i���D�9Y����W��@��	�-̙,�2����~'h%9�aV�N����R7�5��$$+%�V8�
�?������J�����>Lȯ�z��0����Ͷ����k�7h-f�Z���޸�d2ƻ�𫣇�"'t*�G�N���*����Ç,�ͤC�C ��Ӹ�}�z���BB�:��#�
�w��[~)�@4k�p�+~*���e��ަ>%3��B�lm�D^��dd Pl�IY����.��)x��2K'�.��MTy��Z���01a��|�"�E����F>�1c��.)�W����,k���$eW�MPBoB�D긞����n(��=���@�l���!�^AC#n��yq����о}��5��ڎɅ�L�Ь��!�k��?Z��R����(���:������Qj?N�D���9At^8�%=F�sSq���ig��ˎʑ
�����Xʻ~��F����/���A��fG�G�\����~T�N�� �r]���TZ��5%�ғ�k�����,͠�:󏽡���B'�1H�t��"UZW��M�k�Y�#�D�Q�;�(���d1�Y�i�{��ܳ��	������I���'�J�%Þ�"�d��̊K�K���4�(��k��b�\x	��)֪�feJ�A�ۡM2G�@��̣v"w�i]c�C!xy�����DG#����wpɱ �ƅ�4�I����_�Rl%h��<5 ������u l5�dG��&!89�U��	#W.º��)��k?i9yx2}��e𲉣�Xdt�q����B�}��p:�C�&)�F�&/[�E�Jz��..�Vと��l��I�m����	q���8O���R��ۯ^/�+�z�j�Vmm�S �Z�v�h|�;�XSqtikk��=��j>�F��%M��~ԇ�w[�2T#�h���V��B̺j1W�Z�)f��2���G�+�����ڑ�k��z5�%��;�����s(T@���!G����l&�~^�wҷ�T`RQ�"Y_�c�������P��.*&މ�}E�� �!*JJ^>>���(_��[B���㇝d���Jp�5/��Y�<��}`b�Q�����9R.�ce��8��')w��H�.6<�F���nG�xY�ۑ�g����#(�:l(���pyJ.5\��Q���}��^:��V�~��ŌMt��J�i�
-�`^_��%���]�l��ü>�[ӓ�����%��8"^7�y'�Hƭ��d����;1��:U����iN�d�O\�q�+�(>���~W��R��\��P=��+��#Ó��o�[2�?7L���j�c�?� �����bRgO��/�
�f`��m** 3Y��n:���s�x���;�XmwuFI恒�b0-��)r�W�5��W��H�7�oն�1�fA9��e(W��i���Z���8G��&D��r9)�-�඾~��Tɼ �G}@Q���-�x<=��3ʑ%���CX��o������$%���tMi:���2��i#`�N��Lё6��K��'�Р]�ﰮ��vo�Kq�=v<��6�NM\Ske|�bOͤ�U�$���8� R����+�Y.���j�4��'|`��|�^/>��o�	tQ��	I<�Y��XQb�D<[W?� ��0:�����t
b�M��2r���̒@��A�̵żS�Яƥ� ���j|�㜎Zu0�\���9gtS:+ԁ��@vUY1��]R�npmD��|'��c�+��>ix^��;a���ʖ�M{�}�,0���ы*�s%;
QO��)���Ζ`�����'`�Lע��M4�H2Ϗ\o�zv�#]q�z�[Eql:�ؙ�dq� X[!��(=�4`�PG�&�]��(�k����5}�D�f��������9krx�O�[��.N�\�k� }mj S��WE{���(��a�t/�����	�+1(�Q}�T��<1�YM��v)~��<�n���m��MɎHl�¼�l���8����`nW"�a+���J.�YEr�%Q��9��k�+h>-����[��_)��������L�z]	�niaR��$���<���t1
|O�ح���˭E�����3�#�M�W2*��@���\��z����%�Ƈ�dN�c�{��|�؉D���b�>3V��7����"(V��/Ps�`c6�恩�4��o��a�e�J��oK	�F���Z�7�%Z��X��2 'd��Zbń @�P?'r��A<�����}&��?/7@�+2�Cʓz��+آ�XY���Mzܮ��OɎ�~�Y���>W�~�:������UX��y����~@y�j���,�xP�ٵ�oK'�F�[Jz�}���x�����d%;�hJ/�8�9!i�+1�������*0������^(�Foi�U��D����31�f�6�7�ɽNM�8W�[��0K�V0{l���G�fo�Pz��A���.)! �g�3���vDfj��"!������x�tWT�ݽ�'�Hc��"���k�)|M>���0�R��d�U�bؤu�d��E����C`����vWE����UY\�ƹ�>[F���N ձ��5بݴ����UW��<���RdM<������'���߲ת*%b�Iy�PR�`�%����$i����|e���_o��蟞�'�Nx������8�A�@����"p f
||�ώf)����1+kXv�!�� �L�>��2|�B9�D���a�m3�!$�͸R�d���jSGvP��R0.=+W�11)D3�
�}�a��=%�LJ���ĹEe\�8�с�/
��L-�[x0���Y�e*��+�D�.�61�+�/㰞�>�; I�wk�^�5����ٚ�X�Z�2$�2����lZ�#(���'0��*`����D�y��k�6�
9W�wbg �� R��<#zH"u�l���U��ep%f%��Wg)QQ���B������x�����X��P4�)����ז�1e��6����Kb�|*�3!�l��I��CG"шn��c3
t5hJ��y���!�]M\���!^
���RQ�L��"�3�z�<v�f��3�,�
�Eۺ�q�7��_ٿ'�K��D�ڀ�4tF��F�9�"M���ԡ���LE�_��;���n0XʳG�y��3����GS����ݏ�4���1�a.Nv�찵;�k�g'aZNG�'9�҄SPdmKn2+��G�$�R"�ǆ�6�ӓpD`�	�~��I!6z��)J̍��qb�TUO%L|C��ef�f.��
�55H��(yWX�&3��9��{<_���ӅXsdMOkIp�C�
����|�tY�?a�m�%J1w�x�}� ��~'�#���S�����9��l7Q|���)�={�4�'�L�����R-�Z�Q�u�lDY���fC�a�2����S������K�ؠ;!u/BWI%���r�&šy�:�P��Q~��?����Bv�%���3[�L�Z�Ƽ��V��Z
���ęm�Cnx����3Z} 
M���ɕn�J�ΣА[N�
���Ʌ'�j�͠ń,׎�s���,���s;�j/ �>���	\q)�=mSXx��%�C��"�x}X��:8�G�eY��Aꨁh����dD��~һ�0q'�bE����;X���\;��Tx=�xio�2f�HďP0��nO,�����;c)%����Ć@�Ku�0J��D��8��})�Y�[��T^�	���5�~l�͋�̾>�.:!^4d��5=P ��� ���.:8��0˔����N<�^Ǳ�.��w�D Ean��ӗ`M�y���Ŗ�闡ʓ�YֿQי��m�{٢M9�<TʾNC���츩H�/8\�]�<A(�_;1@�3�5�<�AS!��Ǒ ��|L������Y���Zy�$z����O�� ���l)f����\N-�y�ݻ��(�JM�n��.���<��h�т/�H\2�/2)5��(L�!K����H1�x0���M�&���� ��!ryi4���p<��oj;��y��6��/�̮z�c�<���l�D��xﮔ����x��,jݠHI���m�f�]������Z|CgTUHK�aN���p"F1isgBH#Epq:��}��i.~�X��ۆ���D�m��
�uxDYP�^c�vbׇn����2�O��Ux�mDwO]���9�Bt�M��T4������zu%����������	?���
��Y~�����n�̦�mU��qfT� u������u�s'��2��_����s����xؼ�V&�;x0]���^��_�`:���1�G�7�FE2��>�]3�Fc�۴W�D��z�ÙZ��6ri?�*a��G�_�� j@�����gw$~���"�]�(˶=d����R:8k�IqT���V�vggg��Ài](3&d��T5em�
��R���T���y�s؁��M�)��N����I������Q
�4u���4���#U6h���Ծʭ҅Y��j/�X�2�Qֱ{��2,us6��^91K|ob��������U�U����'8�xt�Mr�J.��I�4%�#9�j�!hA6ees�����j��L*ӷ*�q`o�0�yJ��`�%Q����q��Ykj�1������dM�_םx��Z�vt.c�'�C3����X60�[S�#�A�$/�tV���̵���х5��I�oe��6�3!~W�-�O-��k��WH�trҾ<�Rʾ|�F-k~v�!�ɒ?�*�u�� �P��K�* B��#��׵9W��B�c�֖8��ӗn��[�2]AO�B���Cg��}m��R)بk�9	�A�VSd���LOD�P�h��������1[Hv��f�aDD�-�ҽY(�?3'  ���v���^}�����I�(��'��B�RD�/�O>{�~%-eV������_���w*}��b�釹(�py�����q[��H=���_\\5߅BI�,�}<��4"#�������s׶f!D���ttR�q�?I���Y��Ν;�-�|��K�R0(D�'X�֖;��!��n�$6��yb�`�?a��E5?X!��Ù���΍�-�3��e�%����Xn���(���z����D�+�������a���@���t�u��lf]�g'&tP�E&2x�=�QbX}�fhɄ$ᛸ14�^���`�-��h�����I{Z_�C.�m.�u�q?�t��3�Δ�~v���OG �S����S�G-vE�?5�9����偿҄L�̶B�1y?�3C�MY6��-���cՌLrxD�x�)�L��\^W��x�לϰ�e�f�ʊ�� ���6%x^��宯]k%��/��Q�o�ΐ/�ͫ�Ĉ�l,⧰椹݈�	q��V�s�I�fD�H��(���,ٓ��@�uI)+K��<�{@^]ⷜ�+�hr'��0B�YAh��9���sU斎�Η���'�.N�y{z�g.����1~E6+��g�5aA�4x�B�-��&�DM����4?�ޟ��x��x�e�P/�-�{�=�����+�.���ûCjS�/�ɕEg|���i&;�{�7Dt�uq#�n�Wy�?RU^q�P��<�L�w�N$1)yk�߬���spp����Vi(K��)�DXfn2P-��S?�F�����z-�ƙI�z0��ڠȚ<ƕ�J��������?z����_�keHm�LLL�g���W�������~�M�E�EK�
��3��[�[ݿ ��:��E�<��V�;��+ݻ{i��Z����������Eb�2_H&+~��dFݼgҾ̭Wx[���j���d`��o���� ����I�'�џLJ���oP�W� P	�Q�M7���>;zgZ��?L0�w�Bf O�/9)e�2��U��*�+X6o 닋ж��]�9e*Vӏ�ͱ˘��E���OlQ��>;g�4��2-δ}�_�r���5�o"]��ŭ�G���7}G_I���Y�-]7�!)��
@55p��7LFL�m�	d��II��[�����0���S�b��*Y�;[x����s��X���x�&|l���񷵵]
�6�n�h}7y��+��fhO���AZc]����y�����=8Z���P�S��T���_̑q�wm9�VcӚR�>%�[1Q�Է����7=�U͟��[�*����(�(��D��	�=�(�K����-�!V�w�w!���Q<���1����.�d-H=E#��{�0Ң�M�(ɨ�Er8!�����J�zZY�ܷ�*�~h���� �y��*h��ts�!D�VԱ-/߾��|��t�O��ݳĖ��
�Gئ&1᷶�zή��$bKj��XG��c$O��9݉Z2����\�VVݑ����M5��"��c�p,�B7έ8T�\	}�\}0��q��g$ʥזy������d�)�N ����@	bܣ��`BZ����Q�3ꅁ�M{K	6��(D����y^���2'R��6�p�k��F ~h��%�:%1��/4���3���f�cfηz�r�}HM݄N�_\8|*��K��"=,�����5X�?#� �}3T�p�_4!��<��*���t��>l{�q-�c�{\җ\������4�9H'5�ҫeV�T���h��wk��Z����0Xؠ|6�@T{5I���^�^l��v�6nx�s1.>�gd��.�i,��DI!���l:��bBB��)�MڃcdMoư�F4�(<���_��e�%����SR!�9TR�hq��D<N����c���62|�� �x������TB���IV�#_��ߛ���M�toF0�\ޢ�C�Cr2#&v���2�i�x�o$S,�蹺FN��Z�&c}�?��i���g�2�\W?>]t�Zg�i��3r���x�ˋ���|�����|G�����W�݈J�5��	��Q��}�3�	`�jo>nۍ��P���F����ռW�Ϗ3�t�xZ�¼� 洸7\�(�۷���	��w�U.���4$̥���]�%�@��̚r�\�gz'�a,��8wB���+��/K�Q���Z>�P(������O[d���N0��OP�Si�li��wtG��y���܎S��ǒ��l�Ks�:��Q�Wd?�8�0��s����TtI�+(t���#�7ؗ�I����\L�*DO�����S��,=�N7~+EG��qg���b��2}��39[�eLXzhQ��|H��乸/0I�j��3��4b���L�qF�R�x8ĹAJ�dImÓ>/�&�QK�F��jI���(�B�/�	o�(t���3�P���O:
�-JF�w�2�6*Jz�l��r[I����-:a� �cN�_�7����HCvd��꬀�Z�y�,�"�Ad|V��}����c���D���oI�+����!duoz�z"SM�gr��&�i�6�G��{AB?�ð>ksD�1�9E���;LV�a�.{2��T�.'�|q���~+�Z=N..3kk�Nӻrrr/�g��Ԁ��A�`Zt�S�R��������e��^V�h���b�#��|_�/�N��?x_��o��&^����f<^��L|g�1����&�@̞����t��4�1REǘ�DM���]K5�y��*��4Jн�]ylHǰvk"�=�Kt��]��]?Mx�\��P���N��ࡄ������N��~��7%%i��2���9[VH���J�]��HK�ʹ�ԟ��Q�ˆ�Z����|�.5�����Res~j�$�x�%ؘ=��͵������<<�_�W�$`�U'|��C�0k,�H9Nq{�PG�k��6=��<�:����5b8�N���1~S�f0��LNFi���}�ק�� /�-����½���jy�Ʉ��ʤ�͋x��D��!F�*U���$�:�h��oSih%��|rr26�3s�1�>(���t�0�g�t��g8K��D���?~{ϛ8�qx�����i=�����y$��[x{ {{6�8���un�~��}����7�X.'s�	��}q1��_�.C��=1M�Ľ������x�΋f�vG�:[l��ݤ�F��)�=���<�����G�7�/���k�v�Uq�U?�:����W����^����5i�^}�D��%0��,����K�5ھS9B Du�m�`,��?ec�ޙ?Wʠ!���E�<K�5��l?����>K�!u�K���VW�O׆�}��v�L�^���u:���ɼG�d(�%�o�u�=ǒr	�KW���,@�raƹq+i$�/;��`J��N�%�
�[�����oc,���}:���g��B3��wf+���L"0
xݘG,����ב��+fZ��� l�%Z��9���Z<V)��P����)b2�涠��nc�Is�
+g��'�o� 2�������r2�����aee%\}�A�i��EmxV���u-Q`���Q*���U����IM��K�.���|�B�d<��Ԃ�(p^h�	쐇�ƫo|Zg\����X�0�o����ӾI�$"����zq�$u��v��#|(���;�X
eLV3��_�<2��6O�9�4]��Z�L����n���;��xeܐHu��xa�X,@ս�K��휲/��{7�ǒh�*��ڦ;虚gb�Ix���o�q..�uHB�rO��R�L#��Q��]���rU��*[��ek��8�##}6��9�Ԕ�ش��VP��_��_�[0Rx����CY�a#�A�&S���U��D�U�i�P{��g�n����M�^�Y�����<�w�i���x~t#u�?�CN���d�����Z���Oj���*��+�Љ���
���1��{=��ּ��9��VyS;�=)�lB��GUC5_���������ʼfV��gE� ��\n�K;��"���L`��)�=d[����9�ܭY
,�exu���<�{�n^�\��<&���*�$�h�������?�3�zw^�8��I)1taXB��t/���T,�j
W��B�N�L�ޘeq�ȁ�alK�������/�v�>/Ϋ��B���f>3�&��^�,$?�`����x��2������v�#���,O��"l�J74nݫ<ih#x�1�������z��w˲���E��Qς��^��/��2�m1~��̊F���È]g?���ۯܒ9H�{G�#�J��|��F���Q��-S+T,Z�2)�2.�WO0����r\؈'�� ����2��g���;��x�^%:$���m\�!���ʖ}��9�o�u�s~deQ����F.�����ڐ������Ͻ<�)ꙿ?Vܜή�$O�$� '&+湓A��D5n��V7�y6��.� 6�skf�cv������R�˿+���j޾�^y�df��B�}�7qV_l�R��D<�s�S�X��JPĮl;��qՂ[��Si�=JkkU)���1@;��X罚դ����k��t`�u@tHB��J1��Q�u0���@	��(�:�7n�K��^-{�ɹx|qִ)��	؏&�1Go!��#���T���5��;�^T�W���L"ӝ��!��dxǙB��@5%EC&���O���IbԸ��|1�G�=`;���+�D�隣T�p�s���Գ�I�����;���[#-�:C|�M-=ޡj<1�yy�
�Ȗ�1bw.𥪡n����n��P��<��������b�t��9��5e����"���/�ˀ�Ve:�D(�<�{��K�J���p[�O��u1�p|�K���J��떈�e��֏���'��q���������v��t�wGI��4O�`'](�:k�q��й��9;6:������#������5�:�d��6d�X��ß �$78Q���m�k���e�����s��X��G��	�2�VT]�����9�*���z��ɒ�>�~sm��X�=��q]�3kQ����%���t��e�o�K�G���FWaX���MԜ[��
�2��8&?_�~{!JOa �����ត�go���g�FĮM�~��Ѻ�����lɛ/�8��Z�n��Kb��ީ��`���`a1��ᩚ�kJ�n��G1� ,�]#l���Հ5�f�D����"�~�[G��&����G��Y����n˗^�[�!��77"*�I���!%���l�%'t?���b��d�FEw&0��.�\{�e0�E�"\�9!'���"��KD���^����_��?��4wooAn�D��xf{D�����ͿJ�w�	�L�"���MR�0���N�9�/d��u��Q�m��DLa������;Df/}��G&� b9� _C�?��F#�q;�=���#�:=V�K���c_����1�������%�nr�+uo-�z��đ%I&����1�B��yoX�X�n�>�� 1�UB������c�'T���7�o�0]n)�W��W�nZVȗ|0���4o���r�oz6vD��H�����&O�������ԭX�2tT�k҂�;:�x�6q�l��8�䂘�;}�%Hgև0A��ջ������L���[�zDIL���[��bS3k\�M���F��4����x�)0�C�l�Zч����8!�Q"�醠	�@��뿩��r�i�A����"2��'���E�/��p�qݸ���݈���� ���#�o{ta�����Y!���v�C�f�_�<p���)򬘓e_��ޅh������5z̰�� �:?�g _�hh�����B��X�=��>���6r_'�HǓ���u-�J�=YT�C��7ɣ����n���ݜ������ׯϊ����e�]!�=�5͎W5�K2"��/�%��9^u���;�~+B`���#`Pj���r)<��\�����"�3+��J����.�P�sm�"�珹�����k4��{���qr�p�:ȱ��<��oG�P($4�:��]��:c���H����>�r(��H�7�̔����;��s 	[)d���<���Ĵk�[ގQ�|��$���pk�1��W+o���k�{�nё{_�{Z��?}-93�zu�B����ER�ʲ����3���kQ9���0�oN�����������x�Ƙ�-r������۵vPy�i.�B���w���2���5�g}k�� v�%6WSS1�( k�(v�|3rs�4�5�������^㠿��{�^�����vǢ��A�ǟ�;�y��f΢H֠� ���#�F&�=�[��l��}e˯c����\��FN��O�[�����M�v8j	����K	O&�l�| ��3+���H�������ż�/�&��p�x�4���L�}nn���}�Sf���Z< ��܆E�!� �!!!�����r��|�oa���V�є�}�u���q(�
��Sf~-�N�p,g��0���ew�#��=�$ީ4���/���J�@h����Ѩ�����$,[{VK>���=M��MR11�h�3����oI�H]>��4��&�җ�PB:�T�E=L=3��}��ЇkFW��=n�a��	���~Y�U�gV
��p<*�L7����.��4�@�=�����%4m�^���]�/��j�@��ok<u�+����FN�.�WBp��QF������gij����d�J|	��W'�����^]E�%,!��m�kr�ezV*���덑O�H8�|�J�Nվ	����;###j'���n�(�8ÕX6����%����n�3@��ތ��U�Ă�z�_�ѷ���I��u*����t&֮�Hn���Y&j��?�z��Fn�%pK,}����)�*�	��O^��q�-f��y��!2��]�\�@� �X_�';��.ĳt�'G����kg�QoHޱ��jr���S,0�40��)�᜝*��#�p<���:��Df.^����\�o�%�3ry���宧i��1�B�M�|Zv�h����ENn�\Cn�y"a�Z®^�C�;1y�Us��u��P��Ml8��l�+2�+���\*͸�I�7�́Y;�P�����PW5?��j��":�aI��hoUI�%��	��烜�����fݺ�u�"4>�=T�R���~��;W�S����\���T�ً��j*�o#����]I��Z�峪��/B"��}���"�A�V@�K7��a|�0n��8�:�Hrb�R�+��>�0�X'�֜�Ϧ�ż�<��-��V�<2��SNQ��9B]����ӞZl"Lv��rˍ��7�	�s'�v0��%44��M�tq����۷ؿ��w<��,9�X����<6.:c_��	��w�ۆ[�K�޾�'�}u�H�v����֋�������I���*�<oL�(�nѪ^�߸���Ak�R"�EI����F�Qx8.-%+::>�L�YG=���d��6~�-#���~���7#kv?(ڙ�p�B��"��d�Ԙu/mp*����n���.^�whG�����S��GSx���s�����G�#[3�
����X���w��+Tx����+�G���Ş�[�����Գ+���$T	[��=?ښ��<#���#�8�]t$�.��a�գ��(��sK[YYy��a�B�px�cll�]r�^���``��N���[�6�Q*�g��P?`��*4��6 &_��z�P��'gZ�{*�;Hld��z�彇���n;ɕ�͙FD���O���-U�Z����P�ڴ�JV�8a88�s��i3�^��hȧ�A�<V+)-a�j��2@V;-�/^���#�2��3����C�rC�[>KY�H�jsq>�8�m�i� \����ɚ/^X<R��|+��}���c����P�/>��$�P<>��k����'S�SQ&"#��������G7/�����˽)��`d+m�Qn��5O~~�=1/��sssN�����F�.��(�`�?�jI���QQ}s�IN������+��B�6�Uk�*('�Ɵ�+�H�!�������q	;G]3�����ޥ#_�f�۫���m�#n�̈Љ���a��6��:F.��׷�[�V3ic��C98JW\��Ց���Ę���@��||0��d���w�*'~u��=x𠨼8��>�<C�ޡ���IJ�����Kf7�o���^�4^	oe�q�����$٣K�K�CC�No�&*��	O�K�%���$��۽���ldD���wD>|(1��C��tތ�إ��J���&6���ZX`��Ĝ>�.�,-�����="��yf�w�
Z��㽣.�0�t���>O��=���>tq��Ue�5��n��,HQQ��#�	�T���'��t��v~_�7JHH��B��VZ#�H����#�;/f���s�"{CP�_��,���^}�͘��q�?�-��n��~:�Ǎ��}i����{�&y���ק/��d���f��~|���m�sy�-	!��.���;��r\%P;7=q_��y��/
�Ca�^�S���kI��&Q��L������C\֝��s7��N:�&ߌ����.�G��Ĺs����[�������t-�x�M�"���Ցi`u���7�HII9%~���굽n,L�ܴ���;� ���yH������S�jռGCNxj�j��+����)����Eee�����GsV�;�����������s7�<��zs�ULҧ��͇a�jjD��]������_��r� ��42rB���?�9'/�UG�^�ʍ�t�+���	r. ��.<�A�D=Wh+o��?\(��Z�H��Ŭs�
��������^w���uҁ��'E�Ȁp'//! 	$����e�pj�����������b�b:�+'��Fx�ԁ�Vp@M����_ˢ��?��K8}ݡ�~-I��߿�7qr��ǁv%�r�w8�i*7��>PMM͈;J��5�}�[㿕W>$��	�O1�f�T��aG����ÛH`��%��2�����py*���j�l��*of�W��,muu*C�aCQ���Mu����xLKۇ��N�[}�D;�+*bS�}�i��Z,FH]�������q�*@J剚���?�5��T0�I5�M���^���O�ޭ�v��=+n�`��c�z��b�g}��>i���#~���[�&M2����]7_/�{_�l��z8�ω��ɗ�4�ץ�zQ�^�Nvf�W�׌��k�p�N�*��-)�����+A��xr�	{���w}�%��.^�F����[������ ���x���^�A;��W�GԻVD=�KK�s���o+qb�׳��N��'�g���;C��'2�wi��u��3ڻO����*��U��VN��,��������#��+ģ��������]J�T���Z�2w��D����ǥ�|�OG����"Wo�p}Z��?�)q8�=���D�χ��������f���Y��Pm��R���HC�xгT^Pz�F�M�(deaD��oF�3Vb�O�^-ϧ^�嶵{���h�����I��t��y��������K�\x�ׯ��iR�{r�g�d���Q�(��7C33����������<]uXU[ӧA�)%�A$��tw��tw����t+)�]"  ���������>�W��kϚ�Ŭ9lNۅ7 2�a�u#*��:��z��0��'�\�/^0	��hY�;��5�pO��#5ൺ<ٞ�`�ۗ��ln��I�ic_�9���,��a`9؄��׋�<��!���H�H�v A�##��e��M���X:����e�[��{�`^��Ȉw==R�,:*����L0�^i�W��b�_�oAUU���}�}��Ľ0�lF�(X])�+G��@�;�քu�=���zv�"�us2i��mAw2�$��l��BGPS�7y���|P�yC��[�ؘ����֏�z.(��u�$t1㾛��֬�	p%\���ttl�/(v��e��3v�����+~=����k/o)�x�)A�G����@�ɯ:N�ƉN�ы�]]�@5m�޿��]��ݜ������M��,���,�i�=����3��Қ��O�j�0=3S3���;��fb��~y��jM#=�_�00��)�����'+��ܹ��2�������A9!Kޞ�2��&�����[UU�vrw��f)٥yi_�B�c8�� ���"��ĵ���|`�b��W5Cr
LFt*V���^�<S�:oG�<t�F�ƣ�J�@qF���N�oP����5r}XWǯ�2�Y��l���Ň��]��?�q���k"�~��32�B�j�T���+=LR�0��oɜ>����������f��U����j�QHt�(1����ܲ��>0:��F!i޷7����qF;S^���m5��}`�KM�y����d��%���`]q��#�Z�2�J��e(��<[����9��߿���C�?b�x88. �I��V_c���\�;����d���o�o�rY�nf��c޺�L}��u�O�=�툤�p����2����� 2�ꏗ����q����E�������D����_��.��t���u���-\�1���
�L��,Ȃ�@�Q��é\��,Z�f�O�����lַ�sk�����������QS�ǚ���LLKիɥ)�^]1��/�֣�k���˨=�r�M}U�K&��o~T��̛�zG��:����O&�^�_B_� �I]��<8<�q6��#R/���\!O,�crd7��Fۛ��I~����,9
)ܥ��Å �	�>VN�(���Qsފ���A
��8�ؿ��0��n��y��4a��ͩ��xNƌ&I�����닋�u��ۂI�7�s���2;z�`0����гt���?=��ҽ�}�H���m��P��ɻr׀�\��,�Җ�~��f^)S{? ��޳ǟd���{"9�������֭�6r���ˈ��#��@��Ēf4�ky!#F��^�W������(���,f����{E��+��ǂ�WuF<�Y�>	c����C���m]�d�zt�뺌?eU�Qѽ0X;����l_����I�S�W蒤Ԥ�찈���G�i�+^�냥�)�^��œ�q ���_�~B���=��5�؂<_��,(]VnK�����o�*�յ~Ʃ�we��4`����@�N�_�O1�@v��������W�Qn�/�T&v��ϫ��L6�^�B��~* 0=� ��F��HC�[J{'w̼���������P�m���R�(ϐ����<2�*8�����BN[;1C�]�q�6	��?�љڗWV6�x����s�f�Ad����|a��"����[}O�����ݚ�D1
��ee/�؁����C���ּ�<���^�5�-�JJ�I��jj���&�� ��ݎͺlk�w3+*����s�osf7s���ǉ�����`�n�'Iw쪙(�,wढ�������t}�{_�o⿑p�lmm����H{X���dX�m���&��_Y{_�$pY�$�ki���~[�헒��gdD7��pʁtQ�8��J��2zm�d�ɧܴr�Ҫ��	�hhh�>��������0k��Z�I��$>�_�[I^�L�Д���O�^��܂F*A�j&k��o'("2����5\�&J����a�K��u�dOv�Q߁J�x�L�y��r�#n��D	 �U+��O��=���s33F��2Ҙ��,���E|>��t3��5�g4�E��,��6�n��ɸ%fhH���� ^��h��F.pB�3b��Q ��D��c������^%�eI8�����p��R}��SmҚ[�`�X|R5mE�y��e�~��_n~�W}*�>�����}1�2\�=�٩Z� M���¦�p��}�Hq[��GqF����{���N+=�-��X�x�Y��2_]�g�Q`��~DӞm[{�3��,|�cJa���:V�ˋ��f��hVkn7�Jf�P�[�,�W�,s_֔��@�^�������[4��	}�K�u^�/ �1QQ���&�0�$�v�q:���_zs���-w\]]=N��'I3�N�cA���R��E4@�j�6C[�F}�y�V�����q��C���N��ީ�k����Gp�Okky��6�~���cz p.��ƅ��<�W���V�/O�g="��W;6������0�nMV������d��y�'}4_L����8,O�z�ٯ�k�v�p��|.��i{�6��$�"f��|FU���rs����<�?X�=K��1��\�@1S�C6�?��@��0����cM���������6�ܒ>�Ǐ� ����D�6bH�US��C
kj���NP�J��j]�*^�m_�=�[\���HX������jZ9m� �l�g�� ?��?o!sk���������tֻў��hd =������I�	��ht6K�b\�D�H�!4�D����X:��bz��uX�Ţɡo>O8��ܕ�������V@Pn��&��55��&�ׂ5��:(�����J�"��M�L�8C�̼<�����l!lzE��\��`N��*�`��4]�Pׅ?S�*-�7FϫZ���O<�9S��������r�c���a������ ���
�rc����i۳^�{i��B�*�9zxZ�%$���˟u��K��w�ƶ�Y�α�X[�Li�l�u����IW����^�p���Y������o���A��>�o5����9������ݻ�F��>jj�W��_rq���9�!e0e��rv�s���A�g��	�KRW�n�02�
q���vF��@�.ԙ�* )��w�9�U�zH�����#�k���}�����v�+���҃�ee�KJ^ �P� �-C�OH@���ٕ<t
�:�����V���u�зTc�p\%9�|༪���LP �b��+	�%�^Vd����Of��ā��R�٣G��VV��g�7UOv�s��� Va=��QDV��۹�x�K瞩�Rim��w�I����=��l?TQ332�ɟ�����#K7�|�+�N%��o`;��5^��p��#'Oe� ����;�yJ �P���-)qq}�L|unyl���^G�#�;��k�L�;���nt^T�9���=U}5�{��/#vbb��j�p�`�ʖ
�3t��у���������=��l��{�?<ڱgI��r�@րt�d�/�[�&��U��}av����vd������K�ތ�ɭ���7���.K	@IZMM��ժ���*_R��/AA�ㄨ@�^M�9|̄��M��Xj�m�0�Kpp��0�/�������|觔b|0�z`{hd��v�m�)v����$p)��,;0P�̂ b�<��i�G�;�Ui���-㐕���f�����hx�M���!�������T�3`�� D[�P�����zF�ӳ~0�ˑ;;��$�M�������¨~�7��Dk�EGG�T?�@�]P������� R�a``��W�	//��[i�u����	�����)99�F|s������H||ǿO[ؘ
����Fgu�k>�v�v�n����z/�WU��D}CM�=&��yW7k��z�?b����G	��z��zL�բ^靬 �*6X__���Z����;{.��I�a�-���>f�)7��:�0>&VV���U�'�߈90um8���_<���Bx�h{��k߅? îv:=+K�����*&�vyt����Z'��| �)%A<2���T9�d�$F�{��f�|�*w-...�|̮���̆N�'GA���!��3��u(㼚�zO�գԱ�읉	@�<$�v���;j��v�i��KP��<qt����T���%"�_|nAM�����4���i�cc�d@�����u��'�����WdC�)�c� ���	Xb� Y��lC�Z�ǁ���X5�d����j�J�hʂ$5+k����d��~`c`I�Cm�?Vx�^�֌o�:�]�<���U���v%앓j���Y���$,I_jQ�i�2�nMתD��D���jj��S:������M����z�.	�L�L��&͏ 3G��oQ���n��7'��4c���\\���~X�y-rw\@=x�^ }�<+˭-������aͤ]vvv&�"**��@8�R��UWZDD$+�?�+.���Z��LL
\�i؝� g^�74̀쩩�����-�Y���'mg �s,�1�j��qd�HFϞ߬$X� e�уA����wAnė;ZytD�����!k�z�'vd�����Imy�t{Fp�5�č��7���4 m'��
p��;���$K��.H��]#ʴ���)��cϹ[��1k; �v騩����n|���T�"̥44���6�R�O��%"`RקϬ�Rύ�o�hW<��4���_��<���	v�F�m��xI���uvu<�Y�5取u.�"[�w���F�����QM �f-<�K�~oPL I�_����ΪQ����đ���XЃG)K��g��=�G�W1LV��Z��[�{Dk}FB��������z!$�^m��jO���^ɻ��@��`����cٍ��t06���l� xFx�����
>&.��o�0�B�*�� �{e)�'�q����O��|-��b�yc"P�s�S��K�g�H�zA�>ٕ�����&&���z�;@��o@�4�[����|#�P�(�nY�j22�>-��j0�f�v�b$�Z::X���?�����z��C�J��vt���9�C���]�M�17R��vH�eҿ���<����Y q��2�<@���Gӹ�gĸ�m�w!�ǘ?����i�s�������BxWbW0�.}�Ch�|�US�����Cmj��1I����C���bX�'+,+p�IA�p&8��ϫul;�nm��T7)af,�&���������gʥ�l����^P����Ԣ��t�iv��}or��}� ǂP�~||���N`�����Y�l���0d$��89�������9_�ӭ�p��@�I�nLQ$7P�����.O����P�љ�P{�uV.���+�`-�hj�:=3��L]&��a��;�#y�r��Qs��J<{��Nq�9*�m-tB&j��Z��}z�?�)�;�����s�$yӛ���c��WT�\z��)Yҍ+�6x�q�Gg��B񬭿��3��8�w��
��(x��,����ܨ8��W�0ix���wm���`>�͢ckaҪȻ~d����#3��THr<��k�ۓh
(3�M�̮p#g/H8L����
�ߚ{凢1��s�Fb]d5��N\a8�.��M�_��;����cm
bd���I�S�s$�p�A�8�C]���"�i+n�AD����!�$�����mg�V����.6��}�*mT�I��w����|[MK��F�b١Vy YbX�]/QNQC�(<q��z&�XnkrB��/�����V)����}@���iϙ���m������_� a%����4th*w�]9k7iYY.T����O�� ]--) ��+�-�����X�B�����yR��z	�9$bbbm�ہL.��-�)���@��{�^�Nv�|6�Ʀ����zno��l[��H���h��hS%><2)�O� A'`z�ȸY���Ǐ�ި���R'c!�������i�cB�����?�Y��u}��}s�� ���/��9�T���0�Fׄ%%%,wg7-@�P9W`8,s/�0�.-/���'�����\�z�9۸�E��� ����9������Z/��b=�q��?3	�7)��?��22�>����u���	�i�I	0�d�G��t�z�JDћ�n�iR��۴,r�͍��\�����
�"2�׬�����C������<��U�{oL�[P��2n�r*�/"�ᛶp1���_BC�=�[L-,��Թ�0�·�f(f�!xxxf��ݾ���AD\� 9t���I����U6\���)'�n����ԔvA�B�l#��j�sE��l<�zWS����f"�LD�Bm�׊<�����{U󬸬���u�t*H�:����U�d��.[߷�OZ�Jgn=�<88��,��x����cTV�'W_�컚���4%ܴ��$a��{�~ҍ�:Z�j��W���p��r���oBQZA0\R���^p�}��*��asE>+��$\�6�"���uu�4c7.n��*""��+�և�7@�2�͜��wtw��_����V�:��!��xm�2�Ev�<`W��� ~��~���{T�(D�N��W��MD]C/���ws��&��M4@XRZ� �؁;
�$QN��5�3�6��Ѻ�<fE��](�x�ׂ�Q��x��EEC�v�a�n
j�{�'ݭ�0 ��:��͔&{`N���
��h|����'��*�N���o�\��~1��@d�
b� �r<P+"^^ۼ�{A��	��P[ʥ��گ�Jϟ��(e�p=Xr򋈌������]]��b1h!�6J[o�ܩ��~�
�������<�CJq/M���h�%�z�1[x�9a%<jt�5t3@Z$#�޷Mr!|yUU���+
zzּ���FQ�f_!�w߈�
Ld&���-��VP�ʩ�S�V��'�]Qj��Va]ˆk}i3b��z�����&���3~�G�b��*�������Ʈ�G�hH�z��0��$ɤ����\E�綞��D2b%��P�}�O�}e�uZ;;����b0S��ǊŚ���O�R����?*֔6#\9U�Ȱ/����@���--�d$��ԛ.�7������=8d"-'+�ǲ9�Q�=�*jw�mVm�QF�┨}���J�p��FԟV�.�~��(0�Iw<�?�v�'/���֏�i[Z�ψ�z8f�р���O(��x��?�k]��^u��B��ǩ�E�o�3�z�.%����������7��� .WED�ԇ�Ӎ���A�̘[��ʩ�J�Q[�� �jwkHZ�&�Ճ�u�`!E�u�쮵������%�rLB�����}�M�޴󴌲���\[�|�U}Ml)�O=���ЫPMz�Ӛ��y��R�Ƥ�Ɍץe�m;�7�]P>o���[G��|��5e��^����`F��4��3sH:��tp7��tvJ��{b��l���e�$<gd,�7}�A�뜆J,�o���)]"�젋��w�؍w#�'�1�z���((�E`��M��.�C�'�ް�fbd�ym�������t�����������۷�xx`�I�f��>����.�FiC�˼����e�� ����S�z���`�%H�v����k$=rN�K'��wK>�}� �YMf~�/�o<<S2�Z�����J�J���g֪P�o��&�쀎H:n��+�3
��i�U�l���ߣ���C��bo��q�uZ�����Ǐ������m�$�2�@�+N���B�ۋ�F�^551QQ䜜�
�\4eu�lb W�1Z�<�ĩ� +��b��l�v��J�8E���Q��^�tttL���a�JIQ	L����f��n)��}/�� �����r�� m~���8��:# n�m4܈��c�>�U�Gދy�=e���6{>�����E�9��ڮ�Q�j-@g@���{CKA�y�;�r��>��ח"�V�q�|�a;g�1Bs� ��1��,lt�d��7Q,W���yyKW���{��^W;΍T��ᖗ�-�������L���h�3��[��z�r*���uVbXD�����k��?&��f_Ub")t�6�
�v/W�s$���X�oM���� ީ9d����~D-C�u�RZw:��x������D�B��|5ž�sT=��l!�u��ݢM&��z�(M$`��,��kO���&��`����(�(+�pF�]�gb|x䄄b�5���� 4�h ��-�J�
CSqכz̽h}w-Ul[[�?������� 'k�L��TZкy|Qkgk+�W.�V���I�6Z,���>���/1�V�W~�
���6!bٜ/�L��6�w<DG���3���f�whXXzf�m���5����?�L9'1j1�B���/�Ԙ��~��DY�b�Q���D�LS@p"VV������9���9k�Q�Tv��/�$��rǨ�;���6.�1���&�L�Gkֆ�-�?�R�������s��D�i�_ܚ����m���C�H.��ga���v����r����5�Y�4����$���y����:��������o�����y��/�$Mfo&2�PͿ2�Q�9F�4K����q��9��Ñ	�c�ɟSP�rgzW�c��_�l/0*�/�SQ�N���Έ�{U�4]dj<�����)������o�Bo*B=#ѕ�>_<���(����ږPqi������'��4^ �!�Dq����2
�GZ�/4��z|��O�����.�\���]k=#�^�Nh����:������J��W�N�ù���i�?b	Uu0_�����=N�1�P�_U,`;���c3M/���F�A~�[D���C6,����
٫g�F)��]c2P��Y 񛬓95�����(ЩejG��iyT��FR!�n�ҚB��J�Mʹ�=�*�`���PRI
�`�݈��t̙�m������݄��� V�#/�t�>���W	)�M32��~;�`���>\FF��T��S�� ]�9����7����"�L畟ۭ���,TF 555�~������J�Zq{(E�j�w4��H?����2j�����q?i���.�Gv�,m�N[RΙ;:w��,@- �tt䠅vuRٸ܌JQ����&s���v�a�����E���+��t�k���1
��(��?tx�u�M��ȥ߰��MlIN��g��^F�O�����@H�}�_�RL>�q�A�.̍&�?���"u�bˆ�&kk����m��:��W1�A~����q�> K��c))�E9�\�se�@[:�kj��������j�# h��GʕSa��:��_&�5,��ߝ�}6VdP5mՅ\L4�^ϝ�)T+Խ���p�}��Qa9	M'��D=&"�w'>#�.���>W�b7;C_ұ5�����z��������X"��t�}"X�.�������������Y�����5�'Ww�gl@�W�\�~���$��M*%�����:=d��Jw�UXz:5$a_	u]|����| oh$�bascc��]0�W�>��>"��G"�ޠ�U����b�k���E��.�:w ����ٯ���%����YokFA>�������#�������ռ�k��e7��C>[Ug�Gz�ã=�o͢�d/��n��4�(���R_�4)�,��P��V�04��^�F��[>4�������}R���u�W@��O�"E1m4��m�u�Ӹ{ӄH��gَdl��/�_���=��L%� �v훚�z��`��\UWW��M&P��f!�U-�!�"؝�����N����51�Y��ۊ:�] �@��u�B�㽱/Mq�*,�I'��n�څȯ��'+,f����D���K ��6p�d�I�i�!��^�^��c�j�}�_l����&m	��c`����	p��}����+�(��@\�lQKk皮v��n�'���Ĥ��j�?j�A�Z��}�>��#�Iy�BM7��e��?�<�l~��	��wu��q"������S0х!������ݷ�_��1����-��j��H�3�`�βF����Yn�<� [���!p�% ��pt=�Ȃ���n�5��H�F�f95����^��1SV�X�{O�6�0w��IIb�y��x�����e�F�R�����f��ߕ���W����K�YXvl���g:���-��"#�7sh���m�����q��Ā͊!�͜��gt��o�C'�k�MLL�����8��v�mh#�o��յ��7=�E���I���#֎,���K�<��r�y�?~:�,x��"6*���z�E//A ��A���yyy�����u�#Z5��v���R_����6�\2�6:��k`��[���T@���帑tPV�2�o#[6eS?�g�)��;{��X7^W��m�|��T�y����aaMF�TϞ�U��Wd{�v����t��?���\X�C �ڿ`S}<��k
!�� ��Y]���l�]j�*�E�q����lz�O�>����F������H����+n�5��ci�:��v� 5WRR�d�,~F�B�͡v7�U�!�����Pf�(e�q�;�3�Y��=+�NR4�H_8���ZnN�+�a��w?�w=��߿ԩ��!� -�	y{%����A�7tp�)H
0��������#��V:1�&|�IS�Ӿ���_�x�!�����l�%��D=~1
ϗ��$yE�Z{��!�H�n����\���q���P �/�{2�1�j�e��DN�ʠȠ�� �	SaTC�q��kF���|z�Dsp��Gs��t(���r���&�ia���- ��RP��O��4$Ua5��WHh�jQ��)?���@��z2�c��$&u!֯���>t���ܬ�+���ˮ>���x��-q���P���ϱB��i���'&4���>��I�����:wx�f���l4
����1��ACEETYY9K��pUYUu���:X��i���4��C`ՃK��N,��R�k᝭2M���~����v���t��`N0�wt䄆�@�
.�|"�����9boog��7����k�� �b�UM���m���a��*Vpq�F6�X�С��ɐ���1�ݻ�#Dh��}�-�`��HT���+ ��<��CF)�M4�ϟ7YJ�<�ef���B_F*����kn]����� P��<��$X^�7�t���X��<ٻ��;�ߞpҥxD��� ����o��DGO�Pd�R^ZԹl�3�q�ۂg�z�,\ �T�sD�k�A��c �
;8�4�БJ��(����(^jzz��L����X��	L
�t,�/�ݗ��-|||������RR�w��]��ky2�wg�+N��>3����x��F#��(���/yyg�ף����Mc�a��Φ��&��#eJ�X�:��O��&U$+�����;�蓒�5�"W��A��q�3�%L7Ρw�{$��
�3:UU$�j�����G1�Nh~����;��oD�$%%��M`5^� ��;t�_����̱_ţ���
�P�J�Y��y~�a�ԯ��#��eQ勊D�)�ؔŘA�E���G�>[��_������|��S���~�b���P炞��x���N#�+����W�q��;t�� ᒞ�l��*�m�L�K4v�{�^q�l��w��0ѿ�s�NE�lG4�vP�5s+���m������R��z� ���*������ѫ7|�ZY�����,�u�}�F�Hr�f&���q��#�I�w���׮�������L�%{GPdqqq ��䕕��n��X�жs����NV/6>���&}�=o�L�g�{]�� ٚ�QPV���3:P���d�� (98<��خ/���%~��1P}�Y��c�ά0�-�G@1��Ovyg��?���Ի>PK�̼�� ��൫��C��W[9�(�<J+����s)���\�՞����N��~`�#""���bI���� 󯠠�7]�r`���}̣���R ƀP`��^�R8�sv�pB=��4� .�'S��8���0
֭F\l��m����aG��@uR��eI�Zș�1 ������m jh����/�����mП
� ș����%Y���� y��]����@(���s�R��l��h��.�F�g���-Q�G4.B�Э��ˍ�)�b��k�ww\��҅���:�l����03�������266�SyanW�M�tm�A�@>� ���>�b� �s��P�d�!l~��V�o�a� �(pg"Կ���0�uE�9��8�"8��uhh(,2R���5�wz [�'�j���Il22�.V�$�����?���!�77�]=��\���OĂM&r`@�dg�d����c�<LRԡJl�ς���Q�T�+�W�'�{zP��.���͜Cd �k쨞�t������rs��V[�������FFFP��(XP�C���^y--)##���`�,JJ��g�
Ą4�״u,��&����
hF�� T��)�ҿ�t�y��W9冞�q��%WDL�������;V���edx��]G���V&�τ�(
��w6� V�&~��y��Q���9�ql����9h��k�<>𣸂kaK��S����.r��^�|�<ldò]k0y2y��U����Eqy(�͜p;��"�!�9�
�d\\�%����o�6
��߼ѷ�2,z��*��(yC���_����9ڙN���gV��=Ą�;�����J�ؘKi}��䵬��@��&0� �|��f;��^f� $��\F����Y��x��ѝ>��4�fa	�Kq9��Σ�����#��&�bH���}�*tH��@����[��CC�DY������:s��%w�{v���,�t������~�MBWd�m�FÝ*J�'�A��C	~���uIC���w�ȦZ{�rEP�g�S��k쩖1�.��1zPn�wy���Vw��ش��fa	�5c�������ⶵ��cZJJL?�U���,/M�;� <��PK�0�O=Q"�ũs��+�f�1z�%jbB��m0��*�����A�k��|�}'`��m��ei�&�0Ar��3�
2��_`��7��,��c�jCm���Ђ�
�	�oCtX�ס���ڜ��w�!d�jj/�b�Z��(�-g2��d��F��3�>��hB	P�`�����$��N���i<��"�Y����W �)��Aj'��06�HQQQ\NNh)��n�3+55UD���Z@@�������PK��Ҳ�i�eoΛLR�w�C�n�X�?�g�;5�,�W{"�fz�A@-�����upp��(��7-�8�rtt�W��p���J��ͨ��_���q�6�����Ϫ��	]��e�e0D����\^^��ÓWU�Y��fA�$���{y�p�VS<�.W_�D�a� ��k��D��^^�����w���$X��2��ͥgbz7��	�O@��xɷo�gx�خχ�y�!x�m7��U�4�F�){OL�{FЈ�քxs���EV���I)���\*P@ K���	.���'��)�o0��bS;��kH-���]s�{�|c�����b�\�=�;C_�N�FUն����۫��ď����*�5�/�#�n���(�klr��Da��u���;6ejCh�b$!�Fޗ�lqQcg��j�����99-��^�|Y�bd����ݠW?�i���gHzz:pi�UU��yԊ��1!���Q*�hhh�4j>�kU�ũdYN�����E�U�846��4��@,�o8��Eݗ��ֻ=-��zB�O}�P�@�C�~���AܒS}�`P�U�Te�/UW>W9��]�=��dT��,��S��d��>�( �!!��ོ	o!B�)9�hHY�9�q�q=��tU2�+�\Zf>��H�U�`�ג��p�F��6��D���Ү��P6�shm0�oǇ�K7G�~�ZY��p�22�n	%&�j�}x�"�]G�#�DDz��d��.��`�m��M��6�O�}�g�1O���M/�dz^�`Wo����U�w�\�y0��������-AM���tп�}Z��F�g��IE��b�M�=C�y���4�v��[�����eb��6<���pq6�=}h S�l�d�U�Õn�<���N�(j	ū����A���j=B��f6��	1Opeڥ�����ާ.���z�LǺ̚aQQ�/■Q����)�g�T�5U�����Ufr�%"h����v}�G�I?%VВ4���>cf�-���lY�Ni�Q+��^&&&��kL>�q]�)5f 6Q�I�3u�;d7�Z�W�$]vg>e�D��5�q>Q߱��9�����.�XÉ騯�G6��4�>`'p[g�U��s=\)���z��>^�h>�8ժA��b6^B�K'�<j�r;����'*X���"~�п�ɥ��Ǯ(?��4++�	��RKW�5N�{�N�SV�$p���������I	�]}���Z):�����h�;>CS��_*��=㦶�n@�B�0$ᲀ�x��`�����͒%�q��$����P�r��9x�V�j��]���e���\�aʎz)w8�z7��DwL
�3���Q?~P
^n���p�:mO,-/+��3lI�P*�����D�Ԥ[��T���aE��OA�j�����=���=ի{ͨo�Gu�j���<���2�b��|E���4P�j�+6������}U�	�ّ#��3��'��j�/Rs_Qv�A���T��"��h����\����.7�������%��#���84C5�CZMJ��W�^��;ߜ�b�.�=���{���Ǭ�E��m��v���Nb�vT�OA'�]�E �9?$��t?�Q8?N��3Y��֙��nI'���\z8^'�����Ӕ�懾Tx�]Үp1r�� bV�@h@�T��Fu�*�U�����1�[D��$:������v����N��y,�ەӲ��F[�ni�E�zT:��eU�:���UN�_t8��/�
�(��(���r=�A�C��SH����NXM{�Q���̻�W:��s�ԙr�#���o9#�>��z�sns�3��DX�K����[�����b�Y1�(���xv���>�U�1h�.�x��S��(�#U�t>'+y!޼0-;���[(Q㠱������3t@���v(ڌ����grp��ծvooXz��;>����7�r{���Q\�.�~T(��ᗷ��|PՄNʉ��sYMhA%^�1��.�=�&E�S����Տ
j��4�g������L�K�� �h�6U��uu�&/u��5�b���Z`hͳz%S Ή����Y� �7~wE_���������xc)a�3���N
��^��|-�jP�O�W�	��Mo�\�����-���%����懩*v �r�^הR��׷�P��O�,��5;�FZBd�2���
�c[�쓂�"�L�PW��f���jU(��lOFZ��Q֔��6�:������᜴�OS{����|^̲?d�^���ؖx���'j	��c��-�1`�
�fa���t�8�sV�W�yA���d����,0PQ�1�4~�GDI��ĵa�WT
$A�hE�C^�N ��YΧi *ޅ�[CCR�˽<zrM����.��\~��T�Kx3�9O������	ܫZ֋�~���޺v��$��4ۜ�_�j\�}�|>g|���Ϝ���O�ɒM�z�) J���뼶)@%��X��>��	�,;?�����-b�0#���F:�������A�.�-��ր�����i깡��D��T�`�3��p�y�;&��T��}�>Wٔ�7>�<�
�����yH瓳7m*F����iA�H���u,76�]�ng�g�c�I�P2j�۱��h�l�W�|V-�%��̖Bo��0���Lz�ȿd3��8Rs��$��
'��g$�5�F'd�ji1�n�ɿ'lU��
�E��M�O
|!(7�g 6��h`u���������z��'u�p��r�ڂ�����x�&�Qt�%<_� �D �u��4̬vM0?�mb���OBe&�K�A�^��z�sh�W��sT�%S�j�,H�����{�\}:&��'�"�-]R_X���ub\�g���OCX�>�`���N����&D�.�D(�A��9.X5�r�������Ĵ���,|������0I�;���4|�� ���Q����?8/uMq��o��L�)��3ǎ�\�أ�!ɗ���)�O�(��s�ݕ����Tp�k�t�	�n���gG�����H��~�Rx4��-y��U`�f>�[���"X;a,���b�����B�$%����\:�QI�6�n�a�E-%�@��t���e�0wWZ�ԯhR�J�޳���7!~�N��L��6��k󔤤�=����j��16�8>G��'R/�%���T�N�4I�4V�!��j0���Y��^~{��H���5���<�}_��mؐ��6�����F���J�Ke#N��/�&��N���BXcF��0�~��`�k���Ѳ���Y��#^��o߾�L@iz}��޴��_�т�l�G�B:x�Ѓ�	���.�PcPp�^�z�j�v�[z	*�Dh�H:9��%	WH<<}��栃ξ��P��i{H*H2���K6'=X��IXR���@`���,���d�g�j��4 �a���u}2�ۮ-|[���w�Ys�R�Q���X��VW�Iz๬g�}���4���zVWuw��k�.��N��%\��(S��(�U�Ua>�8s }Ax��Ԇ˭g�K�S�[&+��OM/V�ʸa*����kd'W��4s1>�S��k��4���~�]�
���z}���x������($��Y�������l�wYWc�B����=T�u$�Wp�3������l0����vH��)�e4��RP)\�Z0ay?�����Y
������������iL�+�	����C7qS��duu�[zH���e��.��Ύ-l��R��8d��@�E�1�n�@JĨ�S0WԴA�1�3K�c�T�����g�0���q��7�D^ �,����
������fg�B�΃�;�g׀'�!^ǔ�E)w�(�j��$�Z�'Z�V̹@7C#5P>���ۂj�_G[��u��bN}Y)�d$Yl�4��qL"�*�	��%�Ѭ��U������w�m�
e��^��i�r�J�]y=��(�BW��'�i>����-��Yb�U�s��2���)����E����H��|@�/7��O�'�&p�2�شn�dx�U�q�-��[a9{���6-����d�y��%hp�k�Z���Vׁw�Z�`)�𻾻gʫ�W1�&�(S�m��[�7e����6޴.��.q���B|������Cq�'�͹� ��K�w�2"f���_���ǡ�h��w#y�
����RT"�I�����8�@��x7��9]��{I� �zl�gv��1�f��+�}t)K#�V��R�M���B��z���_{_����=cƖ%ɚ=cK��-�Ƅ���|l�}��K�	��Lv�d�l�G"dɾ�,�������y����o�׼�^�}�s������s_�>�FA���_}Ť��1U��}ً�V�	]y��9�rn�B0ܡ��"���^��&I�����ϰ�	r����<�>�"wP���f�h9Ǟ��\��� �vuBB0�1�Y�9U�k?{�ڪG���^�-�O\����=���9:�����>���^�����An�U,��5���p��w�պ���'g|E��e>I.~:����x�p9����!��7���2L��'�ᩥ���s����ഉഋf�"*�ZX��?x�B��峓]�88nN�rP�������@Y���\t;K!����ݢإ7g8����_J
�I�ٕs���~������̯��l��
�Ƈ���%}vO|���X��l�4W.6I�hO��k,���E�*�ە��QTNK�9��1E��O�юг� ��E�����I�E�3�8�ܺJsH`C�``<e{i;Z��Z�x !�3d�ƦˁI.7)�p�cض�������%p�kp�U�����\
��*�Mv�ū���/���Ґ>Z�qٛ�Z4�H"9���3E����	��V=��(�\�LM�=�.��3�����Ժ�of*F����n99޸E�S	���1} 4E�I���[k��YX�šL6=����+avNP'��˕ӗ~4����h6
���:d��vn2t����mP������}�n�;��������~0������>M���ӷj�.I7�5mx�����B�N�V^�e�2k�N.�U�ER�X�$�-����f�j��rt�o2��O�DZ��4.������m�:�.,-m��MR=9�V�\8�2Q#�j���^�+����܃k�Vڠ�I�6y]���'h���ŭ���^y������L�L>��[�bL5r�ZWd�!WB#�������P�c����	�[P���^�ͪ�=н��l���3ŭOIz佖�,F�U݁i�\܊�5+��&h��[X\�d����`��H�JP"�_ID�F �jb�31��n���}+<�ƀ�O�4"�v�

����؉08by�A���k����_N�Bq)y
��hP��P�2&��p����F�[�����_��ӂ܁�
-���5_���gu'Q��n����(@�oob���7魺�[Z���vE����\uC�X�|0R~;[>�1'8ub�C�a�э(�Yt2�A�0���_���E�4f�/H�+dH��0+X��B�/:$]���y������`�����A�P������]���L��#p=��9�b�p�wW��/��?�F�"�ѳ x�|@a���Z�����}����%�K���� �7�ti0]�:����!�����|y��@�E@��:t��m 1}m���V����e]�<��Qo�&%�j��AX��d�3�?$dff�;Ja�����K��������-G��Xe��/F�e��MǑa�HF�fq);;�/�����8�ii�6��H ]*t-�<�ɮ��ydڦ�M�Rl�px�͡W��������&�?���$[vvu�|z$쿓xKB\|��	 ��AA@�L�!� �v^`�Ri{^[�-�R�����0좬�ZޟnT�C�|�!����50F���p,����L�ņ%[D�\ziA�mc�p_�hZ��N�lQ��"���p��rn�yg=B�jY��.$���f]���S=�]"ў���J�S�3 -,yĶ/����M/�����:7� 
�*�r�-O��SE�z eĀ#�����$���5�mq��2�0����dilq�)��@	1�h�^L�-���:�<�s�$��.����^N��YIF�FT�DTm��U##��EO��<�R��~����+,բ�����c>���6��G�K���g�cB9p�s���2���t|��ݕ'@rAG�ǫ��(*j�6�͊������
n�%s8(�c07y�6t3!oz5��n�Z5)�% �Wx��gN]Ǩ�����?��i��.���,����"�!Ҟ	�ݨI"�f���22���o��x�B��J�����l+�Ұ�'��{�QB�ȕ�Zup|=8}Ӧ,��\@�AP|{E�m!�2v~N]���.�������z�8�0��4�������#���`8���tՍ�Y�	��֭q�&���zV zzA��c9P*^�>Ev�z3�Zh����|&W��2֩�H;�م���+� b����C�Cۇ~�qP���ȫ���s�ܑ��~D[]�{k����)	̵cH4d���"�������Q�A���H���h0���r<EH�����o�Z��@- �<;|���NWy�=t��pLwh�r<fK�Z㦿V\KM�u�>�i�=�vf7�'Q�r)W,����]3z�s�l(�p�E=���]b�v c���ӥ�54V�m��(X��3U`�~��!
�(i�a�3>a��9߬Δ�չ��7��H��a��/�O_z����r<�i%��<�V(R�\(2N�o�ʣ�b��wxp7@�-��RR��f����i�޿}��~���$��cPO�Y�)�����t��N�O��P�����I����yŧ*�_0����}1� !8�����@�.fK@��|/`�/���~�Х�w��M����H:�$����s_¤�.4]'�#}{l����ܫ*`��H��Up�Ӟ��t��/ϲ�c�"� U���Ϳmc�N`�OS��.���������;A0��z�d���Z!�l
؜�����=K]�6u_�11QZ���gY1�MI���8K�e���ѯ��R�tPuaa�a��h~��p(��=EA�^�vK�Гo��X�+�|@�W;�I�����G�
٩үZ��a� J�����@djvj庮�ONZ��-YDe)�){��n/0�����!�����QAwY{܅I3�c�A�*����%�I�W������::
��h�i�2ف��5�{�`�6CD��b'[v{�M6t\�8R�=$<�y]�2�z�Ҧ�+�4��{�2�؂�gysWXWu�z�� ��!�)�:�oԭl�dC��?�R�M[!���
iq�`ླྀ���s�d��~�u�*?�Օh8��Z���l����.GD%��I6��P��վT�a�A8���`�	���F�S�@����Ia��V�Y\�"W���g�m鹙�`�ڴ>+O����N2�dۯ9ӋfU��!"X�\@�3e�H�s� a���bC�{4��o�@pD���1d��b�z��SSS���ύw�m���El� �/�Z�(v����Cxw��	�ba'#B��G�2���C���9��FO�D��7�4L�՘E��A�6z.�䦆��^�l+#��j���x��]�Q�A
Z��P(�c�Т��d�T����V?E�c��p��x�b
3o�Jn��:PY3��+�L��ôM�y��ɷ�;��ב�GCN�9z�gu��M�"�	�g���^=iN�ru� ��v�Ս~4����פ�.��pwm�d�o��Gz u���2���`j�QI�g��8��6��V:dmuAT�{!&_j^+M�)�4f�������b�e�jL�ial}��vQ�}0��!�?�(�gaV��{�|^�B��wT�mIS��(Z�蠕����
=�O�#V�n���s�-4�%���r�<9��i�V{�F8��vOk�Dڗ�����wɋ�.��|�xS���h�_���U/3���_Ш��Z����E�LX��"�pND$�2��6���ԕC��E�~�菞�1�� ��C��8�4#�LH�t��V��Q<�X��zԚ�LJX	.R�ZH�w�v�v&���x�O}	څ�O�w�ec�6��5���`v6fr~~��pZ�%�U/����©s�Ր�5{����#��j��@i/�zx��H���񢏎�1G�6��|�$"��]ow|��x�kC�K}�f�
IҪ����'���5ގ J`̛Ncu��Ĩ7]'j��}�Q���N�v�rh�� ��p[4oOh��~^�P7k��@�'pMm�\	��t��f�vܑ�;�W�W�|~є�g�2.e^s�J�+�Zh�K�]��4Ew����W~؃�E<M|���F��6ºu+~"	�;/��! C�3�73��!蔹���
�]��cj�
ZO�N������|�TIc�J@<!;}�$!�� 1+��p���Q���R�JA��L.��>ƨz�$��6�D��"�k��5��O7��(��'�M�UŞ�	W���2Q�>�Y�����R	<�� �%����f �&��˅�_��VC*�ؚs]ޯ�k=U�m��)>dG�(ˠ�)_�)�Ͱݵ�E��O�MWX�����f��W����t��9C�n�X�̔�JO��'L������w'`f��n|�[�*Ny��Y��b8Ր/���[�1:`o�+(r:I�:�+B9�=�}ȟ�,F�HI�'~Zdfv��U]X ��P���2��P�qAKC2(����S7�����)v�] :@�������?\�>�8:x-FC�&1{i=)�>0[���~փ���� �0��k�R��G�Y�gto�����vJ���
�t�ƍo-�\����gN��L�(6�-e�?X�)���2��Z�Y+�1���RS�;���dY?��J�)))76���?Í�-���$+�?��M�b�%��C���w�n���A�Մ�+E�J��m��2���쫓C���J"����
�e��D�dL��!}���>�ޝ�m�-�	m!�nEsoܤ�Qt+p��o/�j�D��c��iy�:p6�Ɖ�J�I�X��o��W�H-�*��?HEy��8��y*",�Y�_�sOW���l׏��G�_�Z�1-U�@��rv�����g#W�5Ѫ��׺�?s��Alӧ�eq�Q���ڄq ��6�4�t48���=|ǋI�J^c��sF(����b�{C���T�0��2>��@��݊�<��8 �nS��H���R�T� }�x`$sf�b����%�P_�Q��%����-ܴ�<�t�(�X�-ƇE�vvv��P4��>~���J1����h�4�Jk��)Rt ����J^���Ԡ�3J1(u�Y���r��RS���=� ������Y~�sY~3s�O�CJ�ź q�nS�߫y@*�Ag�ా��ɺu�ޒ���� Nb�A�_ݰ��e�-EQ���`R���$]'!9���&��<
.�m��/6��; �o�����R3��P˝�o��j^�V��7w��ϐ1B�Dki�:ɑ�[���`���jM�r�t��.���߾W�� �_- y8���G 6�c���Ҡ���V͍�[h%��f(����󹪀j^noQB���U��.�H���C[  �"��gKR�9���2Q�g�9�ش~���
����wh%¾�ϯ�m � �67��7;��6����hK����^5�R_����ۤ�UΪ�՟��9�*�o�5���Q)��FDc���Z%�}��m B�o�tN~��u0�5�h����8B?���r��7�f�.A5zr����b��C��EO�6!1�]�^-����P�
X�I�'v `6Ж�}��6�>ӎh��2|f��N���d����͏�8Ж=b9A�b�m6��|�=����+m��A�p9>�{��  ��Zw�f>Ȍ��ZP�Tf~J��Yes�wy;�F�	��T�Ԥ�pZd-�2�v��;�q�������A�e?�l|և9��
�)�#��Yч&wk�+��B�*��B�ʃ��#�{��� P����M�㺛��k١�C��!��IIg�،t�$XTOj��#���?�!�b���ݾw�����jP�߹�ɂ������-���r��y9��_0K֏8u�o��kMS�����B7k7�=���C	�����Io�pD�jE[C1W�?{�E�j� ��߀��v4.�85��*��Y�}�h�E�0�)i���ŭ��4]%!eV%�8:o�Ҵ�N��H����Y���SyY
@��)'L�������c7nz�>��:Hn�C%�bbљ��� jmL7��g�5m
������XjQG����h��I�b��7� �9>�3�9aPE>�,`���n>�?�O����k��(�G��KWt���.���'<>,��Qr�A� �i'	Jc!M��p;%�	Y�����ʗ�)Ö��pL�}���O�u|-�:��6U����dd�h7�R�ʨ���qp�9�^a�g37b�	~v��k�z{������G��.��mQL�����d����Jc=ah�O	����<�,DT�*ɺ4�߉sN-�G�4��5���*3�����7Pp����xvٽ�XZa^���6�b30x��ƍPǫ����g<_>��W=��f��}��]3+����Ӫk[YY��"���3��2sb\��p!(v���J��V�Pspx���F���X* n���S�ډ�<zs3t����h����'�<��GȆ� _������[�ƴ<Ƚ��������$��tC>I�%u�ֹzbpɠqp�ZD(g�w����]�}U�e�k��3P���o��m�uI"q�E�8$�N&�Ӧ��g�uS��0�ȴ��PW,C|�<w����U7�m��eIq�I�� t`՜9j���]�Z���V�X.��yG�i�@���@��!!��L��CΈgafl��>�C�B�w��5�#bħ�]iǵ��x��L�(*�W�'Ǚ�[�u��1�~���
�h�����r�]eL����>�BȪc6�G�Ŵ�6����j���K� -}�@�t�3ԝk��QJ@a	(��i��-�%��^����?$p8���/��}�d������ ����o���AR�	w�Jj�|��H��|�Z�(����FQ��qY��W���q��x\=-�R�؆�{���n`��@���q��/���*Ը�p[�xk�m�����`���%p}���bL=z�����u[cB���7�	P+�]���[�Wn԰�IL}8~�h���S���cp����=���l��[ׄ��]��d�	�R�UL�����Y����K�7N��oJ/A�p�߼Y��&P��6�U� �2�|�.d�u���u���ۏ8�/�b�K�zz�P���>�������ҷ�]��<�t���bt�����l;>��+J���c1c:R^�h�~��h�������0�[S��g�o���<���ƥ���~���l���Y��TQT=�I$e.O�P��.}āp��ա"���ɴ�,ȥ��!�`��=|�l�i���ߠ -�SPY�!�40��2���{�҃�LS��4�jg<cϳ���L�1��L4؏�ǐ�̬���?���c���O7)��ur!G�����p��SVuX�����lt1�r��$]�w���M�R��_��H�<��(t^R���o�]�{+�NV�`��@����.t�|�m�L�#����2�%f��J�qr����)�WQ�m��Ȃ�e3v��52�M˄,������)��
��\WX����[���6J�t���U�HA.pՎ�de�+���i��<U�&�pf�HtFfil���3Q�;�%�)Oa֫el�k*���|��iĬ�[���DM�L�����1��e����������װ�6��ƬCz�(�-D���$�&���G��u(���RNhH��0j��Ʈ������E�6Z1��������*�z�dhst��O�o�1���ueA��*i�9�H*��zpM��24���=:�9Y��BՋ�>M�ض�M��h�oȦY���|���m��nX��+���z�e3q����{���u��PK   �rZP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   �rZF���?� Q� /   images/f590943e-678c-44eb-a174-3243ba5f3820.pngl|	<Tk���ܴ*�})�F)�2�t�d�2�L������'�m�si,Y��kBc�Pѐe�C��4&��4���ֽ��}���u�s��[����9�~�і��!��sdS%"�^��I�J�<��}���z�߽�7���7x��BC ����V5:_6(�ex����������__�C�n(��u�C�w�Rg�d!��c�?/��}Ƥ�X�P�#�}�`bVO-NX>��)��l��T�z?Jo���c�!P����[zl����e�Kyĥ��j�������v(~9�9�D�FWo5�`�~NA�L�L�4�M���-;:�6RT��!f�Y� "��!ɱ�����?�snRr�D��n:��8���0Y�T�Ip��Ҝ�Q�A�-f.u<��}��Ha9�:�C#J?~��X��s&�D�W��t|�ljt�X�g���x<�K_�C�LV�},�2�����Yw�揹ճ�<	WF�x��C4[K�9�p��8�愝���c������4r�3�v�R����X����i`O���-��LȊ���G��	H������hhiu�r�ׯ_37lےlY���~�Z4d�6�I�革��)%�ͩ�Q�[MF�)�OV��n0��X3<S�/}K�M�8hD�2Ϟ��s������ ����~G
+���i�j�[ZZ�c�cta���{ZJ֡.�����m��cɵG?�Zpm���k�����9ׯ>q��U�X�Y�P���Y����_P5��a*���z�$LT偽��;4Hè�<H�(�?�t2��s��;f�9w�O!U7��b�+]�){1K� ��"[]�c�d�z�0Oa�[����s�>���2(�|�z��[�?�����
K�9n���&�J�����Q:���rrrF�
�^�0y���ݾ��P�8�is/3���CE\b�m�7��'���%젡A�֝��)n�;o$�)Y�?cd4�����ǲ�W���4�+���H�V8J�&55�iek��	-iӥ��PW��*��CCz~�G_7Źn�s�_w��G�m��ϋ~�U�dkih�KjC�]1� ̈W��0�펻�Mx��������$M���-L���{�����u�B>�~�Z��"T�>11�+�������В��8���B����l�C�:4���y�;�W�$#<�$�����S�z~�"2i>5v���Є����� =���h�[߄ɓQ(��	�o}��*Q�=�9�"�V���� �*�6�^�V��k����:LY�Pc31�qP,�«�gZ�����V�vЈ��$�1؂�|�]4z�`'�mB�w�F=��[vo��0�����\�����@������m�W����ю�g|S���q��f?��p��5 3C�_��+�'�R�?���Y�S����GLE�����	Ӡw��qa�d..�\�z;�m�:==m�����4)g*�*1�d�a��������'�-F\�	[����;����k����!�,l|t��b^�z�����*��+[w�ҕ��Slg����	c���or����Z�$�*
��@�����mq��jPG��5 ������K��}��v��q�X�=a7Ƀ���g���C�>k�Mi[������z���$���wk�Υ䌔�|�����Q��w���9S�z
79�8W��7�<����ٗ�fh7kM���0��X�>���3҂�<�B)��֋ZK��uF>&�<�2-hjjZ�|��T����-�2���!�xF���K4즕O8:&|Yp���S�{j�2���t�J�0�'���5�ZwX>��_�/P��3;t7��co�ȉ�Ŝ1��C#T��I��N-����k(�KR�
�:y�q��9�N!�.?���s� ��j��L�b9��&����?b���*d�C4�ew�nU`$aAE�x�n��2e�J4%!�d�.������8	�MCVBP�!���f�U��#�g)�s�]: ��������chu�u�(#X�R�h��M	�%�Ȭ��HE���J�٤<�,�#��B(Uc�̗mo�r!(��	�'�s��I���`��BBQ�K�[GS�dՍ�
(�C�ְ�n��m�n;4�JZ���|٢��i�]V"�':��-�����|K�s@��'��` ٿ�A�k
��~��^
+[RJ*���c� ks�vxpQL�� ����&��4"��Lb�%���	��w�`��i�r��
��"S����-hw�5
��B� �x��՘�b薞��;�(_8�\z��z7 �\����u];#�U#�ΊYY���Oꅄ]�������N�n�.]�!k�ϤZY3�@X��ϰ*9�	���Z9%wd-��m�C[;�Vi	��gR9��YX��1AŘr2�k����I�e�oL�c�c X�� �$��I�-Q��3��`8	YP�UsA��O/o�)hn��]����H��y�H*沠���G�F�'�b�U�<HýN��z�{y�ʕ�/kk���.U�iC��N�e���lmm�}H:L�W�jF����I��u|�OB�*�%g	\N�m��vL�e�Ӷ��I�A�4�����_L/C�I�h�9F���*56�!�UyO,Uc�P�r&MQ�e��5��s�TM�AAW����w�+=�ב�5�I�>UNva���v���������%:2ק;t�$1yX��w'�7��9dڥ������,��ij���dV��?�*Q�B���`�3~#�	�/�#I5AE=.#�}�W!f'a�9���Y����~w�"(_K���Q��
�
햘��2{ s�M-x�.X���%R�NN`Q��,�Ȭ���%�K�U�xʣ{����o�?|�y���Y���Xe��ή���a�3�P�|:)_�T�8:�<�����%VUa�����ci�������ɒ^��ީHP.��=��WJ�����,w�()��
HWu�c�&d�=Z�ܢ��V���~�
g�HR�����J�u(���5����#Y�*��V����g�����h-�4�͛7�C�x��m��w
����^����~��Et�̉�A�P𷾒�T��״��)~ޚ~�7ԃף�W΂��HU�����\`�ϸ�Z�s:��Y4]p��H���q�o			�Qw���q�� د�`u���O~d��2���hJ}�x_x��V*��xcE�O� m-����f��1��\z�[�a���5~���q��
�~���7W��i͚#?���t[�74|q�ҴO�~--U��~�t@Q�5�5J�^�Ч�%���A�Z\Π2�[l0Ӫ���d�_��ͥ[T?/{�CXy��d:>U�-	l�"[)w�#�Ȕ�4\&�Zv��GJ��>ё�Z94�7�ݯhJ3���$O���m꟡�K�$�Q_��Rą&$�R�U;�$vu*���Sæ�g\,������,G�.����ڵ1�S��T-��K��j�#\�����]-�E?�E��a8��C��N�[1�ND&k��M�R-���ʺ^1� R�\)������oʂF  �W�1Z�����Q쨿i�P N3�S8%a*��L�f_r~V�b�+��^��G�PO[ͬ�W�k^�0��:{�R�^�?�iW��,���&�ciG0h���2N%|K���h4���{>4�Җt��C  �L�u�uu{<p�@1H\�U���_7�V�������A���w #��z�Rw��T�KR,έ3s|f�!I�_ܓO	��֥D�$YY3������41�}��OCכV���I"�a8# �G@���,�~]�:�<Y�f��ے|H��R��a.�Ӽ������TA����MK�u"9i���	CD�W��~>e���_v:�v)4�4"�'%x���CG<[E��������圲�m�»K�=���#�$ǥ`n�?�P�O��K��m���Zch��m�̅}�����U1O�"����8���.�X��/s�>����&���50R���V�ڏI�pR�&�Ӯ�y�Zk|��#U��I!�^x�f�pEo��"�!��P��@�f"ml�&�v�릓"�%��"����JZfv+�AO� ���2�a5^-W�K�C	bѝ'���.����Z�r��/ՏرI�u��&��/Țī�d��s��< x�B~�����I=j��dA#0$����Ǥ���P�)�X3���Q�����i�z��?(�u�9M΀ѩ�@M���j�#!��-��G&�dD��5S!U��s��C�$t̘�i�Q��w�_�����1W2 ��\�V@�3�f鹱R����)A���;���p�L~d��(?��%�Չ����G�6���-���p���sI � IKծ��)�U�a�j�T�{�ek� ��Y�_;t�M�Z�L���i���e3	)]A/�;|��?�P��ى��{2�H����h�n�D�00QK�Lm&w�=��� 2�~N�Z������yMj� ���٢��AX��3�OcY��G��~�F�k6=��k��-E�U1��1�맽�ۀ�ݿ��OSu�A��P����U����IU����s9@y�[X`���۩�`�Iy�x�.���=.�\gu�,u�oo7�7��=H���Q9)��p�jh�XR������)	�(�j��DS�i��:� ���j�㳚��Z�Qů�+���n}{�8顰h�}o�����5�Q��3N�GL.'~=O��*�����@%iFFizfP�>�~ke조�g)�w�7������������r���C�?,��<�:~2f\ic��+fچD��#����m��H69ZQ�Hf���}��5��G���OH#G��g���%�H�U]��SIQn��C&�pg ��D��Y��{-�~�a-��䍞�'!3@N��4 '��%���_�jN�j���D�e�_���Am�z{��LBաm<A�l>��~���w��"*=�v������QU�$2�(��cƟ�u���wg�bT��ӧ�����1�9������ 0I>�����ם���������6������3��ez��G[,����ݛ�x����q�׾(�U�[�ܡg��?M),�*�7���L�q>�c|��N���j��@ ������㒒�'%?�H|VX\�:=�2)���Jm��>��=c�w���G�4Z%�w��'�(���F��6X��M�θE=��3�M�E�ȯ�=���j��e�V�1jpn����8^��a"�Ls`7M��Z�#y��?;�~ÚS��`���*�� ._+�R��PL#�yY���JJ�~�c�����csW}�6:�� �]�*���B�Aw�E?}�o�� �Z_\W��q$�w�B�˹��n�F�Q���a
]�����։�F����WQv�9�HU�������/UT�u�LN��C�9W��%��\5_��TSY��>�/�� `^��5�wSԞ-�_�W�%Ri�vĴK���7��P�=������4�J��zr��c�E�ȇ�_ذ�/,������&D|r����^U����o�t-�-�)Y���u-�w�s[�Aީ�`�㼈Gx��م\�;f�\�3��L������ٷ���?�1��ia��y禕�0��
@�pn����Yl@��&Oyvzr�ZDV�#R��f�*��1�w���j�!r�"W+q(:A���eV@Qk-�[������.�u���$�7m4���_�1݁"�P����y�a�Zdem�7I���n�³)Z��2���4_e
	�sN�m�^�.�CjjCW�nm��+�}�h5��N�j[���凢���	a���ǫ,m���K�� ��IG�y�J c�4^E�T��ӪV{_8/�H�7:�Ǡ�<��᰷�#孩\]y��4jd7f[KI^������=ԡk�g:V������s��R��{�,�D�c�����g4�n�X�k�,B��DI�[1��,h�����D�T�נZ�2%����9��*q�N띌a�
��?��j�nYP�q�h`(3SD�"`�w,,N� QX��{��1A{(��G/m��c�xUPv	MMM����}ʇ�˟J�̎�qJ�e�`w5�p�T)��~�8����[��)��I��h��
��AӮ������[bק_���į7m�d����nN��Ҏ��tƑ�4?��'(���oOÌ����$�i^�V;Zf�>?br�'o��gB�3��'� +�]����K0)+%z황*��*Uc�$�2��i��]�I��,Ѵ#����V��F�����SD`�t5�i���ԡΌ9c�#�7�幖A��QOTtƙ�5NQ�J�9si �ʀy��Th� x9����t�aGQUj�Y���/�:H��� Ĥ|W!4"�TUᥛ��z�e���?�!!�E����30{5W���Si-=n`�ۥ3F�����9QF�{���� �8�NK�>Vk�y����ㇺ0�-ӭ~�bG�$ �:dr�4'� w�m-u����G���4\wg�8����y���>k��x�3�ǃ�@�Ք��q�w�rA��T0~Vt�Qg���6G���(��O�U�����y0!�6�ݧ��e�^�^�2)o~�U��Zм5�4Z����V�����$>:��4V
(��1)� I�H�#L�`��E�Ӈ�ڀ����^�`^aVgU_�OW�*�Jޯ�D�F"��OSo�R�[�Ј�=�v��%|�|��Vh��މ�͖5���¿"o��_$��Q���o�v��!Z7�H��S�/�h�C���G���ju�s<I6;���w�|o?iv���u��T�<m^��_ ,�\�W��f����o��"0�b$g�����6�boP4^+�Zsb�W�^��_� �?�.U��W|n~]ON��?�"&�5��j���<P�����"���K
��,<j��� �(E�aFL����yj�� ��a�C�U�s��x����M���5=3nۈDv�AЖQ��|���K�9�k5��wh!i�z\lu�v:��ȕ��Y?��l,�E��rk��w�1c<�p�T%�@\�&.���J���Ʒ��!=B��^�>=	y��42H_�[���A=���������&�
�Ne�������=��M�.�at�J�+�����q�1�w ��M�� ��y(ߢ�5iJ��М,����p��.�H�	�eC#���	n���,�W����a_8#-,�?\�-�!��U^�o�(��tȄl�������6|�I:�Z�{�b~ާ�-�`���>)CA��~I@�LB��D�������g�d�;v�lK�X���l)b�Ԥ��+`h��A~��$Ŗ����ر>�H E�
��6�8hć��.���0���ݘN�d�Ii�ޥ�cV���U�F�����K�c���E���H�M�m��a�_�}3�۰0(.�C��!�m+��!��X�v����ج�}܈_?�_��$�<���(=w��漟�E�����q�n`N�.-9a��?-�/��Z� ��3����Ɇ�.����駤 �`���U�Ӊ��*Q����%�B��-|"h``�z�h��Ќ	f�x�i�\��ޭ
����ڻ�g�c3��R�L1ݖCKZ��U=.
@�ې�Z�����A��Bb��+|�C���C�KK$
G:��h7�׷x�b0����@�i�nz�v�a[��c��?(��-S �%��(�<! y�$���A�!�����),����] n�~�����?��@V��e����.$���ƨ���Q�3W8`�g����κ�)���`O�Y?T��X KF�`6^˴ ?�v���.&&��+����^��g�ysz�n��Y��E@�2A���2�^��p�>��m*�qNZ�"��k���X�����j�E��5�OYw��U���<��@�M��f�F��Jĕ�5i�f��Cp�-�N!��4Qx%h[��2��V�?@�u�܊�%Qt��_:����=���ZXD���fA\¼���ʀ{�T�T�Ϡ.ֹ�C��}�TQ��ώV専?�=�#�3z�W4��
ű2X����h\��9JkVڡ(�{�Vx�ϊB�Vx�M[�(���x�k�β���e�0��Sk�����y��Yf5���L\�q����Ќ�h����b(���T��
���}�M
��g�+��B5��h8��	�;�q���(��Ո��ۥ{$Vim��3�N7�4	���< �C�!��c����	ߎy��G�OH;Y�3皥�����vwu�� ������8�������ɾ&�ed�<<���Mݴ�@64�"%��+�p�*Q�����6v�g��z���+UcyT�P���z@0��qr������)�P�|�< ����~�a%�l�]�ݟo�:V��D(wu�DK���Q��#�G�D���ߘM�	1Ka:w6��b���٤�VӔ�^K�g�n�0��}�����f3	o R��J�	 :«W^}ά���H�N����b�/raqtŷ�T�\KG'���Kt=�s���>�(�S��h^?��G�5'����@�]�^VU-}��7�~DAf[M�kmںv�g�Ry�����s�IRn�O�a�;"Ǆ���fE��| �@��s���7�&����sQx���� �Q�&�!1������ń�����%�H��Ɩ�}� x���DFY�ҵ�K�
��%��,������ͯ�|Y���\���a~~>��G|�Լ�e`�k%����d^P�*�6!�~���A��n}� ���r���$윙D�3^�n� Y��q�~A+8��#��`9فEXD�1�Pk���p�߰0��k�V;Dn���y�]9_D��x��G[�į�_8�Y@ht�++���s��H�+��yo���k���b2e��.�H���D)9��
��g�����!x��a�-��W! �H;�N�Cn5.�^"g��v�4�A��T�R�lm,�S��ݭo&��s�;��B)+�i1��ouEM�J8�ѿ�c�# �]����p�����cW�����u�"��7%�μ?`2s)�L>�*��=�������R k��ja���� ���{XLLX:}b"����ػʄ����9����ukd6�s�Fgܩ�H����u��/.=w<������������m�H�y�<�wU�OU�>���Xw��B�d����ŽO�*�nҭJ�9[�=����d����O_�'��\O���R���|B���"���=䪄Cn�H�L:�ʈ�v��ѣ�j���B�y�o�(i��Wl���?Y욡���<G����
h�c��Z���I��֦8���@���gzC��u�q j5�Nw�����o��Vhp�O�=�
�D�0�t�hĖo��t'n5A��^�3�)ƙ�Y�[�!����F�oO�tp��@��Y���{����}�^�J��T�s�f��A�w�F>)�
��%ԩx����^�u�����-QWlzKo60x1��\�DL,���ϻ򿳃vӐ�� V�IyWgq[di�e�?�a&zyU��mbJB�)`_i����H�O��tǅ�Һ�w����2ib�X?Xj��!{��U�W�%7�<OG�p�Ϛ�e<qMo &_X^\x��5;��O>b��0����/��m��d��'6�1#'�Y�|!��	��3!�����C�f͎��@���Oޮ��D�{�{! 6+���Kx��o��oh�ZJ6���N���6��~{�L�DV2��)�b�l���tU�����9 ���e���U���.��Pl��'�*���"�'77��V�b���_����m�	��Ժ��!A�l�"���@�7��v�wU��-�?���D�|�	����uğ��f�nB3��Kz���<N��2�f=�i��p	2��B�$��)�б�k�Tp�꟝��ֈ�����s�۫�ܤ�H��,�X�����:���]�����.ܳ��
�����"Z@�9R[^� *f�!ݹYSV�����w�?yb��z�7�wr�Ԑ��>��Gn	=�q���G��o�����>ee���+�M(Ģ�	u�H�_az/�ZG�����2�0}�\�B٧<�!��-��o{���qX�*�h�#_\�q��Rz�3�n7&7���>�+�d�
���;`���W���ߒ��-Y'�|Qػ?�o��_�g�����`M������He]݊����1H<����_bQ��ɒXe�z�:1�^�dg0�V���P��<��}L^T}s��u_�3��Fd����4s:����6JO�v��[OZ1�W&Of�Y[��{���F���~M���m8� � ���f�G�[���ɣ!�aa�nn�Z��jm�1������Cۚx�:͉O�ɛ����G�wj�;���8^�B���b��6��s��f}'�3��b:�(��LU�K>���c�x��)ͻ>wvP*�O�Lh-�~�������P& ��2nFUuJ���ʽ�9�i���ʐ<��Zf6����p��^� ���Y;�h����҈A��l�r���1զ/&i�6��6�?��8Nڠ�}���˩qW�]��J�<H�间{��ɣ��N(|���>���E�ޣ~�?:��;x���o��gk�x��vŌ|��͋.�ة��h��)mFɳ蝯���B����������7^�kK��:S�֪(�2���ܪ�|9���Mi/��?����]tyE��0��2�/e�����M��[_\��{aq������I�z��/�."v�#g�|��\Z��)�+{��ߡ{f��\��q�S��+͉�x��ZS��p����Y7#�r�.���D��� C[^43��_1�ƍ0�����7��iڀ����A�<Ԑ~�r�����ϗ@�AΈF��U�ѩED�z?М0nN. w�{ﮘ��j~��d���s-�*/�H���z�ޡ��ba�_��^��G`K�T-�B����dr)�|�X%d���T��?����3��]V�m�::1팤9����P1��;V
'Q���l7.V��	E뷓0I��Nv�}�sA��ެ3ˣU�O_5N��c�m���[g��=��˷܈��p1�ysr��_��|K��桋(�� ]>{�=������{T���ZE��E�h["�P���wȴ�P�Β>�C|
���5m�=����>5��n�/����Ϊ:�q�m�ʠ��dM.5'�J;�ǧ��y��E�=��_��{��,h�����̢��<i`{R^�.ñ^���f��X\PP��ݡ�]D��Z�V���f��}���v����^56f���.o�mT|t���{m�њR.xqN����}����t(�YV4�,f�C�4���ȇWRUu/M ��| qd��o��cR���icVAL�]�O�8|B�J�6�U�ɲu���\� ����vt��{���_�}>�O�D�G��ʵ��UF���?	���ڡ��-�МwW��D!�������'�1?:�d&��hZ���l&�kw�(�@����=����"ö(�݃��J��9��n	m���G8������S�\�瞙���seu���t�p$O���;m� ��]zܑ�������v�Z��d
�ޭ���-��$�m���0ϏD!�m����	�
_KKˑ}�rO>d�>v�s��٪ sOK^5z97q8Z3�0�"Rg���m�(�x��#�z����	;��_���6�T��Y�t��c��[�&�#�O}�7_RϿ�� ����rƚGI��m]r�m�$K�8���F���N�������"��`�	���cEG��!�5g�l4����O���,D֟(��'\A�Ū��h��,��k,�J&	r�ǎ��� )�&�_��$�\�w�9��t��g���2�˷da1KV�f(�����b�)�姞�#`*���H�e(�����W�>��?�#EG���������5.g]���zR�y���{�G�vV5�7�hX/�s�(�����kH���wke='�<�-�-C�`NH��V���o��O�w�ӌ�7��Q�\.�V�1�KK�k:�!d$� ��F��E�v��[�+r��M/����r���C�{�9�v5������n���%Χ�����L�w�{�����-��l�� �H4�@e��TW.�Y˔�:n>�����t���OٗKBC�Șb���%�t��UU:CCC���Jw�]f8ѪW��η�2'��A��2�Zz^��+�Q�CHB�mY�qѵ�U�f����7#e����i��?����0����V���1��T���OF�77�q�N� #Q�������z4znPlvP���?�z�CAJ�?2�c[8��u^�w�$Eu��������$;�j�:���hek�]��A�F8)��L��&��.f0Y�O�7Lo�1�"W)��-'��+�X��n��7��W��:9��l�v�l�{7����8�ʙ��Znl_ac;������⏒����0�G����,(�	��G,��g=�w1�(�@�`_� �A��wI��������sA��P�H62
���'L>�j��1� F}�Z+��F|���4�9�\��K�3E��O�E��U6�s��yJ6v;�N�~���zl'�����?�EC�	�� T���lI����'��7����O�\:�{�;�� ��g*�Ouv#�	W�,bg+Fh��G�%j��.�~��v�	z=)�}�LN5�g�Dz���y��ӏ6��D�������/.��r&ޙp]t��p�-|JY��q�0~2���,j�m{��n2�,�CM�Q��}�H�oq�od���\�?�����5G�i�8i�+?�:ې8$�8��ԛ��I���j��]&w��0xB"�؝�]&(������{��&]_�p?�S�)K�M�KT3`$�Vf>�[3\ lB������0ޤso;��@�0��:�Lo�Ѩ���c&!�q���|jҋ�S���N}i���Ih�ܳ �T�	*Td����>�6'�Z�V��Z���+Y�/����O�ϢEA�K��"NH@6�ʍ�U��1� ��㩝w1>rM��B�11�?LE�j�Q|�8d�WU�:$��s�	����w�S1��g�3߾��_)K/j�+rv;��,#�K�r�D�Fl��=�9�\d���O8�C��������r� }�uO ߰J����5��c*�P�Ig�j�S�(:��2�����f�O��R0������|red������՘Z�>���MȖ2(�Wߴ�>�x�:Z;lja�{�^�����_���Tp5;H���V��\S���h���I~��/r���r ��y��\��m1<�z��p��!6�|XG��U7WegC o/��D��O�?y<!E~�״gn$�H�? G�������K���EE}�QI�/Z���8����:A-�m�������܃�욒P�Y�ʙ����:appǜW�@O�I3N���B�,���$q�5n���A.m�)�a�gy�U�)I>��ᣟ�CT5H�m|t�j��{ �D�� ������օO����'���I�+�|�ĦDa��j�?^H"f�"��s۱�/�[�J�:G�,lV��T����k�G��ÌH�^*�r���{h���'�^sɞ�Y����4��R���K<s�%��V����$I�O��٧���#��	��%
��؟;?[' lM��Ӧ?)��x[[3�	�Q�u#i:Nwj��]Cic(��a��$*���R��v����A*h�Z�&H�o�$��X5��
��_k�6��`b �I��q����3��؈�{Dܗ����E���=65���)Ȍ����*VY�՜�F2SS�����ݸYU�щ)�>��*��������U~;A�����x��������IV�Q	��U�~�OD�v�$��,V�3>A��KU 3k��d�9��k\�V�Ygxۀ�!����0v�
��� �q���r�OC�.@�� 	���$$)��َVkݮ��]2h��֋�<���E��0�#{4e�:���gᰟ�B��b�V���SƽtIK=���p���M��m�����o���r��a�M��	��Ah�x�Vt���U�͸��z3�,�B=��LE^}�h���^F�iq0� �}��"��0���Ji7���v�H�R���G���׌��F�/,��-3�'`�*s�U��Տ�u*>���)!e��`]��#��d�$����!�F;)}�H	`�!d�*x̠����^��	�ʲ"X����i�jR��/�x�r�����F����=������l�x�A�<uӕ���#MӮ�s�UG���� u��%/(���I��6��T�ͣ��)FF�у��c~z�X=A�>p?�����K�1vg^���N|��]�@�)Ƃ�hl w�R�{���
<���0�y��ۍ����&��n�<�����f����3\؏�����mVe?�n�#,���ī��^�pخ��,^-P���e�oW	��.*�|���T�� ؖ��t�o� 0pb�����3B�2�W!Ig�HC�����D���' ����8�7g�}f]��n�%]��{�"�@�q��� ��7��u�8�Zj������FJ�'ϢY1��*C�n�����nK��Huτ���;y��=�MOѡb����h������}]PR.x����&�GD�\u��d��P?r�Z?��7��;y�4YY��RX���K�BpbŖ��v},=���n��$-�w�A�֧����رM�-t���i"������Ǘ����n��G�)+.�p�������{?����ɵ@W`��\Z{B�{�q1��<��������`���<� R� �V�Q?Bʨm���$���=���ksH�ݬ�����Y�(�Q@�u�Ƈj��{-�tH�Ů��`̈́�E�sJ���ᴹ����h�sJ�;���ww�`W�u�]�X<�'E�r�������0�����{�pa�4�يk�O�X��!����n�PJL
����!�9Gp?1b�[/�v�G�w�n��OF�"8��e#���r�X��7���3��l�a���>�����s�AwRr��t��q??��}.�\i��ܛG8D�}��?�C�j�n���Ir�3��m�����귋�+�f��*]�D w"1d$����U�'p?��P��j�Jg�α�5��H��c��x=���"�ݞ�08�^;�p����v�}E�Z�Jt�K�V/�ra�3�s�@<�A�1�����[�%K���2�@.s%�+Պq���,$/���i�}�ȞE�?5~f!�^sa�׈�I��2�G���� IS�FW0W|1���_��NHM����6�`����)���o�����'YD����\���x�>��T��T�D��=+ۑ�i)9��^ٺ��D�p^c���e�Z�� ��9�KBl���b��l���zf��{��'@����o�}1s���a������s�:bu�<.��MB!�M��!3 �lz������"rb���Бs��ˮ�l�j�&P��_7HKNwIJ&]Zæ6�����_��L��gU��*��3�d�f�Ւ,�����W��+�.�g�	���ql'��4�����RX�3�.�z`�~�A4xk��{;�%� �{�����vB������V�{�g|j�.�����
�w+��9B��OE��/���V��!�_T�q�b�?��>#�ȉ9Yy��A_��͖�EK�Y���L�l�#H^�<I'2�Qt+=���򺺈�b�]�(GEy&0��z�ex����k�.�*`4�j��3�'�c���>����h�:(8%g$9g*�F�,�s��-����{�l�m)m"��x��M�9*5(�r�T1X�����S�{��0��8����D������g�ȭ:��� x��e��Z��0���@��>][�wh����ȴL���ؔ�c�G�	l�$�pTOD]WOk��Q�5�{�=�R�*n_/�6X�V}��"�����}��x�<�s7���_O�bg��E��+��$��	���k(TP��^%�Y�T��P�����y����e�oא;;e���(Z����~���
�8=Ӯz��P%�����Ɖ���!����N޿~Rb�<{�`j�?�k�.%b��f�����2V���7��O��"�p9��EkOo�:El��pN{�d_���G�.�'���rk�4�a�9�+�����Kb}�n���DÚ�:�C��"}��DȪ��S��O���o���>�쯥9@��ٶ�ހ������Zu��$!�m5/�ϐ��O20;���iɾ{ܣ$����G��lv�GrGeUy�6�J�P=�q�r������Hv7�<|J����n^��R��	1��K�ĖR��f�5��Y�=�e��'�x�E	��{ɷb+�o��H��I�TY����.����߈�\J���Y�b!��ҀOt4�����M́�s�ǹ��dw�r{����"�I�iչ����;>+�z��+8��eH�|�Qא�6<ᢑ�asx�����N�NuO�~�"_������)�ҧXL&��W�m&����	ϋ&5�Oq�C��j���.�w1�-��/=qX��}���6����~��e��ߟcW����' �n�sE� ���}�o?�o?�4z=�B.,��ƣ�Ӽ8c*��?-�?�B�����!F�xD{R�(EHZ8	��1�c�lz��{P�O�4�#������4���}x��т��?�s����Z�8�c�So���r/�0�wXW�Q�T��Ru��*i8n���{40Rk�x��_�*��U��_�]�K�:����LP��e�3��m2sɮ�:>
��S���8�H����͐�]#�`R@� �C���=�v��^��~��R
�>�������^
2�1�jv��Y���4�:?�XE+�/���`ȃ�מ(�����>�A�_ >9����z&$���>�%	��n:J��8dP������=��'��S]8띛{������oG8��- �D�4h����N��E�5��7��Ѝ�o��!ϙ��)�`���ڪ6�A��*��1/]�/	�
�~[�K|����N�$q�*XbG���4��C{5�)*��R�E~�W/��I��'�<� ٞ���0	ջ�m�����5P��Sg�)�Z%����o�:,�5%1�7X��9�q����/x�!��r��sw>�5� �@� ���z�Bdf R�[-A����X��ׁS0��%:�rg%]�����9���-��U������ "��Fq㈏�ذ\Ҩ��<bټ��sy= �3bI�pU���C�*]xy>�A]����?��w�15�P^��fWK��/ަ%�`tE��!r�Ԅ%?s|�t�H7�h�11�=,�H�� [m����/����L`T�"��uK����/��>�KZ.9E��Y���2�i�u��}��D�:�v�w�=2� u�p���E�\��PXY�w��}�x���v#��<�-����6~8��!��H` �EYJ��,�$�Q

��/�l�P��
)棨��<��$n��Cey1=�ZLX��V��ˇ��8�jNe}6�b�� �uO,���r'� �8�D�~�)���xT77������x�A	���t�e��4q��x�Z\��<pt���z�\�i�:���������k�#�o�U%�GN��K�7B\/��
`��?����=�8�h^O��?҄Q�9z=F�"#�g�Q���������z�x(���V��$�t�5��)��-�9H��4*5�Ց������SMm�Q-������X���z]w����������~]���z]���tZ.�M0��g�۫�� ����E"����Т�AġFպ�u��6��{��sH�]��F����+��p��L�<:r~m~>������䤢}�¬�����7#��;�e<V�>��hD���:�	r#���8Ht'�$��x��!�t������o�ʕOJH\��mE3�{{S&�ƍ��L�]҈�d����-hq�t��^��{�_�-7?,,�g�]�4$�VP(IwQS�[�+�>�]�k�nb)}���/~.&]�K& �/�l�f�~�r#c�^���@>Xr��it����g�4�3\��M'�xH��P����l�����_�1^~w����*�mF+{��\�@N.b���]5v����V@9�M����#
9�GR$����fD���a��4Ĝ��Gg�?��x�c^4r��%��@A&��a�i᠄�X]�88	�p�Lc�<Q��b	pi
��U�oe��������{y�OJw]D�C fk��zm�Z�>����A�]��}��g�:A1w��Ee����^6B��I�����8���ؿ*YZ����`����E�0Jg��L���J�'0-��ʭ
�-�n-����Ȭq�ԟm7k�cN��u�$�KQ�
W�j��|(+��*�nLw������cb���q��Qp
�3ޮ�Mӎ�ɩ��Fc����������`�S~w���m<~G�n0��,�B!/���ȔLː{\��Dt�q_�%���T7^�<�:Er�	v4����l�	eq~�ʇ�����K�D�,y�,�+[�"��YO�V>�|5�\��x���N�� Ρ�y��{�v�7�i���Ga���ܵVJ�/2��F��W��u�����&�� 
�9�����B}@J�G����!���O��Oz[�/�{���9��s��X��B#�p$�*�v�x�A(
�w֧9��I�������ޮ�Z�,H���<��]y�U!���_�ap�{��b�=�B��֞��a�aM�Z~��i��O����r��6R���E+��K/L�xkoQ{V�a�%b�k3���C���9��|�i�ŝ��Y�hX����N��W>�J���V�t���U���YQ��l��QW��vZx�˹����j�Q��D��)���6����S���vn���Lqbr��������k?��Me@��'Nm�'����R?�v}�_a�W�d��[n���:���	'=���=������U��^g��8�bU�8A�(�ȿ�0��.�WK�ޠWz�_\��v��>�YW�X"�Ѩ������L~�"�J��p-��)�d�"�!{Xc:\?s��yÐa����ǧ�6*>�5����qS-h�ڒ�B�,FW�e��������wc#.0>�<��o�W`jl,^{���%QkM?��vK�!?��H{�q����Tj�p�D�ݎ�{�M��2>��x۞f���&�ˎ����ՅNx�ۚD���$�d��IF��×|���q�R�T�Fc�{�D@cЁ��6�\�6VG��Y���q{VG�z��	s�c��h\E��r����v=�a������b?/�<t�]��-�$���g��POʝ1�ud��u\���+JGV!ҌG�O�����+��ri��z�A���&È�\he(J����Q�h8����1ΏͶ�8����W��6�!�֤�����E����im�UL��}�1Y�N�pk�~�d�ڔ�Oca3��Uh��o}��*&�ܴ��'r�Q�i{�|�ܨ���0 �G�qѕ�c���{C�Y�t���!&�Z"^k�
=�k�f����*F~*�&e3�8��D�y�d?���o��re�K���EeM;G�����,��Z�o���P�c�#h&	#�R~w4�OA� �\d��)��|ъ��+J���/uE��W�V�j�3j|I� �ױ�TL�t�i�����6��Lh��V7H�^���D�z�#a~�8O��RO�
��⅏k��],P$׭(��*ĸ�v�_Ǟe=sƑ'�\�S�>8��W�64���&�f�~�o���x�6`����~aW����o�	�r��"��p06�b��΁<6��N���Z�?�x�H ���籓tؽ�O�Kw��Vso��둗�Ak��3T�rL=h$��)����nN���m��w�����j7|�+�O��A�B���~zg�/����dJ�����BaK ��8����ӥ��	$�[_"LD��E�W!��ςcf��D�`-�i�UL���]OD���Y���9��m���\P����X�L������*�����=~�̙iCF�4�I��f���Z������:���G����Ao��U�ϫ�GMe�n"C�V7��G�_�
��PD��ƒ\�g
�pC�RqX
ڟ�hz�,��C;X8��y^��\��D��,)'YC[�Iw�����ze���S��[n政��u)��<TL?_,���2J!�z�y�� ���Ӗ.Ϻ�,�3��d�	�B��r]+.[�л/�mCB�������<���r|�L>���/��],����`=M_�.��ր������^?��ڹ�` �^2�>h&���q���P�x��g�T|�)vy>)��6$EUwU?�<8r��Ϲ��uف�����^�MYub��)Po��﷙N�o�AK����@��Ӫ�(���.l����%�/��,d���Ki��*�ǣ˙\��'�L2fY���*rҙ���T2�r���Q�t��M%5�+��H]P�Dk�'�ݽ�vJ��>���U'*WP�.����/�'�DL�Mj��)�z���w�]�d�0�X���Mqa`e�ߵ,6��w��MJ�����c����F��YW�S��E�?=��3����麌�Bk=�K�.+���wwe�UOπ�@�?��`M��Fv�4C�����^���o�����e�����6��%m)�E���d��⒔f��}L�ɍ���%	��UM�ؐ��y�y3�@ꒁoI�④r�UZ"��lAhr˔�x�]q@yD.h�@r����Яx�t�X��͏��������LL��N[W*����\he>������0�yd �!q*/9p�o`�����*ab�bBr�?V4Ϝ�M����37fZT�4̦�Ӄ�L��g�]�9��o@��)��zZ���\��R����w�y�h����v$A�x��<M%A���H�H_Wi�#<�z�n�Z��>�^ɸ�!X�'���o�jW�~}r���m��P�4-˛.͏`3��+��L��.]I��q�F��O�uІ˞]~�L�W�H�G�.&�g���Zr�zzeF�Q���ۄn�C���*�2?�<��g�Í����H�%)(�-�C�1�#��E�e8Vzd�^l�5lNo�G�J�26�h4���I԰E�
�lR�xq�Ir�^�Dnr������n�{5g/����SGn4�ZŽo[�_v÷.=8e�c��nu6�"��X���uA�A��"��f��EZze����~4yD#SoBn��wŝ#[��#�*��y�%��Hr�.A���f�\����W-Oו�`���@�9�5)@������(����~h���x�?�9<���'~�!���X�W��M��=Q~�*�=	�(�}�;)=�Y0Q!�?����~W��p�{ދ%�ֳgh�D�C�T9{��nF��Y�fZ��N�fǪX<���2��YC�=��Q̺��r�N���8�t��G�Ȫ,;�[��8�!;�QC���UO\Od�!�n��cAt5�7,���Rӂ��ZW_|�󯤴;��,l"�XiT�͝�Q��J�獮��Ωx��R�М�0"�{�F{�TŒ��qV;Y���hh��vs� ��q��N��E֔��3s�j�6��vz �٦H^�$ǆH�����W�>�X��$�����o!�W�wpQ����ug��K�ckrq��'�����zyO[��?L��r<9���7D;^�t=�5��n���d���lJ��OvͶE,���I�v�&2���U%LJK$-��I��������U��*l�/����篏k:"n ׿H�]�o�\��~e9�M�%hA
�攔��з�i�뷓b��A�qg��u	��awY���('ϔ��v�]�4��/�^C5��Yc=�ˍ��U�U��DC�5)-��B�**ý�h���O1�'�{�!c9��������,�c�)��yO@�Z�&���0�2����.�J4������NCi����Y� �-�^v��,�IvM�ӕ�c�ߐ�)�E�v�ʼ���2�'���Kʎ=�D�P6�mZ_&Z/LcK��6���vM���ZN��.�6ym��\��BV������o�}����;�ci�Ip��Y�n���+,�l��|	�z(��r��|&+������q�w�9�G>֖uس�̠�Y�)�ld��rM��Ӣ|��_��K�ݭ	#g�~�`��N�{��]������]-���{?��К�tK@�6�h�K�9O��U㲗SEO�y+!����z	J��q�R�h���O^C�d��&����c�5��M�?i�r��9�|�5?/�z6?��'�\פ(�ޏ���=�Z4�hqLJӌ;��#�Wu|<W��Co���`u!LpSy�y((u%~ԕ��Y)����" ���eM���r[\�3�B�2b��K�`��t[��`����.5����f����np�+һPD��ۧ�i+K�O�aI����!T�l�,M� h�fC�4_�S��4zWS��N�_C&a�G.o��߼$_��VwS�%��4",���0�c�LB����X�zl^Ŀ})��[�50I[���\�P���~����P&%®V|�)����;�.���;�X6Ò�n��=�����,�4n�U�O@��K�ܸf��C�h�/ٌE,�Q~l��2%��cG@����������x?�A�A�X����2��A��Wӟ����Cs�"?}���~�������H���D!��~�b���%��!u�h¬���؊�d�6�QG�v8��{��;r�d�巑��������썻�OKN^��B-���vUBv6�n���e[FD�eee��p�W���iM[aQ�-_�eQ�W�|Jb\YS���,e�?��.D��422�#��vy�$����k��^�2epy�(YƗ��-�%��\CB&�\��%�mc�;h��4�#��`2��1%���(�Df!��4tM�Y�ocW�n���|}+�U=zT��QP8����N��%,�Ϟ>�P�=Z�����ۗ��p[p���XDpx�Xz~�����΁-��>)��VU�[Uz��I:�~�GȻ�nO[1��M"c|@�"�R��疖��4vD�@�#ig����v�c�����a�E8��S'剸!�GC��MU�ZS�eK*5Ǻ�t�%��d�"0�0��3���*پ�.>]������iHK�Ӌ����u�T��!�k�!Q�j�=E��N2j�P.� 9����@�e��V�p�BL�ړ��

̚t m?�m����1Š��}>���6�.)��ǓǮ��k�y����K�R����D����0�ӛږߙښߙ[�%;VP�����7:���%���w��lVRh�ҹ��2�:qִfgZ�RYO6b�4��+���Xa[y�g��zDO׶��b���j�zudb�^("٢�����\U�;$�c�����y+�ZU���&zjs='|�𱫰K����
����;[���b�+'�������q������	Y���b�	M��??;���k����m=�+ѓ/��*�n���;n<���_�ӦD)..{��c1J��CI_P�Eq>�ۤg$]Z��l�zX�J뒉(A�7w�{Tc(����5&CH�6�m;��P.�#W�M5���/3KG��|�e�a4-���1�P�rZ��K�!���a�����'��"/@��Fr��;*e=�R%�����Ȫ�)J�sl�.�)�ƾ��h8]����k _r��8��yJӗ��W1���q�vR�Ga�5j����Au[I�yפw�q#���`�t:籆|��$�IŻ��|���sy��'���JK�:KL���ƙ��P%a��*H�=�4-�D�DJ�����ճa���5� ��5�Im�G��
�lQY�W�|Ϭ�i]����G���h<*�7����{4ȫ�,��[l��}7�0x������Y��4ׯ��p:��+~�pě��:Фc`�Ԡ�iP�������[�����z���f3~o;�V�$8Mao,��iA�D�ܦ6��Є���e4�ee�I_�%޽�pz?�磻�����K˫��m:�4���'-{)�!���1�H7Aط�R�0�LB�y�f�z7ɗ�rz�a�,$�����Y��=p�Mv��m��[58V�r9�N/_�h�ݸ�~Z�L���4ޓ/q4t����+����e��@�\�C�H>��t�w�AOJ�@� ���X�p|k���ɠ��jd���(J7��l�J.�u�y��	��F�X�� �%��ޞ��U��&O#DKx����V�m���:�O��
iق��,�mC�f�C]J�R	~��QoX�pB~l�$nxVx��Z�)ظ���j�1��c�E�-/���3L�t��q��=��j�������&RH�8�h �}�ʇZ����B5)���:#�/He��dG�&����*�H�X���g�($G���@��E��x�{u�U��8z�{�m�^�����p ������i_ٛ����A>uho�+��I�f��H�c�\Z�m/��%���c�@��~Cȋ̮Pp2�;k�����?x���8��c���
ߞ�ᆓ2ߺ��`����z3�/���+�2D?�����(.����7�=���Y�����^�L���m̶����k�z��_�,�{��g�*��9�X���Uk��޴���x+��D�l<9KJ���Ƽ� �2N^�X����՛���3���DZ)qg 棭�~��d�~V��ƻ��^�R��m�S'�Χd%�U��8�
O8V�NIk8�5]���s���W��\ݖ�I��(ga�
g�v�S<	�ϡ�\�YPꭩ�=�dΠ���r�3���+�m�P����TIҲt!����d��Ҥ�ƠKܳaY ��ǆ�ϑj�:�B�+|��]�ʲ/�F~�BW�	8�1{/-5����j�2]��`?��яyZ*�.�ń2,�_h\���������D�����[N)�lȮ��,���D�@R���ld��i'7���*�W���>��\���à�$u�	�y�#L֦��.�
��`C�L�y�\� c���ͥ�P�W?�FC>���C�"=�J�ٓ�s&�{���(�WR8#�h��O�aj�$��E�K�����`����U��y�a���涁>��8b6�n����0��fI}=��!][����VR��K`�{/ �G0����z���R?��DPg>���*���O�G8*�;��7XɠkWj����0��$s���?�[[�Υ��K�=Bw ��:����G��	�ߋn��J��(m��F���(Ě��l���.Ĥ�{��qM��nx�}$<�7m]����l��D�d<n�oT)_iڂB�cʡ>%�_0��,*���\HVZ�:�'u&��dL���2�������/k�/�p�dT�lJAQW��e��Ӟ����ot��6_��C�j`+|�P�U����C0p��,"�0����ND�P7;���Ko�7�qM:�㟽��y��fa��Jī#JQ��P�]M>b@>���S��xiR��}�t��,A����0#5�՜V�&[r��C޿׸%5��5o��� ���O��f�=��/�8�w��ۍ�Y��ġ,�
1��?�I��x� Q��&)����Ē�L�f�JE^�Fn2��l����i&��E�&?�g)����O�ڥ�|J��o�-�o��gV'Y�5�D��U������~�խP�\��t�X�.O(�G�%��u_�u��ڊ��y:���?S��{��a��Z3ra�ݍ�M��I+���8�K��˰�������� em�S�.�L�&�����,h�M ���޳�/��^���a��Ʉ;��"��[Nz^j����b/���������Di��>A�YDc�y�f��*WCSX�ZI��ɟc���5y:K������;��S�-�n6xe�	����<�%���7}�YL*��>��X�^�P�@�6�8$��t�*�D��CM������ c�HD���k2!�+)m�JW?͖����w��lM����\!�j5��=�RpI������r4��b�%���o�Fn��tZ m�5p��!��x5�e�Gd߹�E)`����=^Vm�B��pz+��5�3��Z� ��ca��O/ 09�;���I��ތ�O��z�&�W�Zq6%C�oGw��:��2YGpV֌k��F
��U�f�AM���m�(���?�^(�|z�W:�t����s�s���E.����7�#֖O�}P�wd�^Y�����,./11% ��Xv�I8���y�߷�"u��`ܘٯg���i��AI_=`�s�
&�&%6�H8�����ᑗf�V<��OOΈ�"����\Me��2�5�q�Z?�J:^�t�H���A �^�+(`��м�G(�&[���/?�ɊLj� Mbƽ�~4�mN��zs�@E8��5������66֫����_�5����( {�G��p�˕�U�U���ǡ��{77-#��u�\�r�������1	����=�~	�|:�k��PRUEg�,���|��g�^gc��Uw0�nt���:.[\��
����bCy�sZ#�\�>�^�i�!�:5A幮)��J������T��������ʲy�=�OĜ���z�"<ח3��r�JMgg1�6\v���pw%Т�=��U��S(VMn�����t��I�wњ6����1���I��Q٪�����~�^�n�Z#�jX�GD{����K��=�hO[�Yxs`�g���:����+��s�9z�	��.Ƕ"Rt%�{�C���J0��M;tEZ���P�A��թb����|e[P��ʠE(b]�i��\ýϻ���y�F�#^'g�QtT6�T��.׏+26 a{=�,ǒ�5���v�ᅵJ̺�Z�|Ü)DB��#
X�ӽ"t%��[j�#�m�G�G��q��5+O������F�:�{&`o����/�C;���Dd
::��R�A�ׯk�(Ĉ�#{��U~k�A>��T��Pdvapo�����
���x�������w���%��7���_|�����ƃ��Ë����3�L�������b5�fQWd��⡖�ɑ��//Gn�F�����_E����ª�/ő�>QڍF��"��ǯ_[,2�rUJC�/u�ӭR��ѭԼX�5��gC]ݨ���l��fm�fGz錖��ƻ^��
7�jkkg�ߡ��k�ϝ��Q�����_^lol���#����6Rh0�m�-�f��-���
1[�"#��S�;i+����9���胦��kH��x�!�-+�X�)~4|����mDͼ�(�<�-�x�J�PoA}������B��~�ʘ�ƈ�)�IvȬ��
�����Mm�I�o���E~
���?!Y��u��k�x��'��ʘ�O�b�7ҽ�j���B��i�
�٨~�IJ�VJGtכ1���EC>��� p��?�q�_��R�2�6����As�x&+d�Ӹ��W D�����k~R�뢤���2�Q�g�����'��XI��t�xv��Hjg~g�bL�a^m��T����:���������H�ېV�v��8Ո�=ţ��jE��X	81mܜ��5��]Q!�$U_I��כ��'Ȝ,�s���zZӸ��Mm�TV�[ٖ5��i�.Y�Ⲟ�∱C:�=���.���;�SD�(�j|��xz�Wh(��Z"��w��>���~��ŝcf���#V�^�h�d��qz�kZ�.����1$o����5ɱCqI����#y�L��#-w2�?��B���՚��/�^������gq���R�K��
T���t�N�z님&Oqz�ŀm(
�!�D7�C>���{�稙�����E�4A`�\�+�u����h�{&f"N~E�54��ڂ��V�ϟ@�"p�Ho(ώ��ZC^�w,�ı��^�_M��D]�^m�e=&(�b����T���q\�'4���Y�Q�ʥE/�m
����+�A@\�>��U�`��]`12�u7���y�y���/�����%Ɗ|�V�}�V���/?�Y���T�k%��`X^�U�n���v
�=��Fವ�t���w5W����D�qC]��
JY�t�Z�;�;	g��[����B
��m�?/(��K^B.���6��)��c��%�ؗ��k}mV�G�L_`�s9fL�MNcCʨ��ID�#\c���z��������6�?���,4~Z���T�,����1R�d�u�Lm�V��)���_Ojץt.T^|Z�z�W���]GQ���I��@e���gb�3�����`ڳ�]^�?o���g��,��>���'c�5� ���&P|��#��&ٛ3��Y��4�)��>����R��Y�2�#c�3Zv�S�
wӴ,�����ia��R�'�� ��5RL�5����'$(�79�c	e�1�G�Z�;jW����:T1YR�u:^S��xq�P�{,�q���Xeޟh���oG/�Vr`3�GZs	�獮9Bs7�u��\7^?��V=#0��.�R8ЇQ�xP��r��AXM��9졷R��� �\��(�C,�����E��=_q鷩ě=����ej�D�2���{oA{�-|o�}��=�|�s�_�X:��*����C1qu�[k)R�v���Hw�3����;)0�q�<��hM��K��
�5&�Ä�|��uwF��A�a	L�B�# ��Ɋ�Β[�ү��!��E�$D���� sw�w�dH.3d��x9�Yw�7�n���QY�Z�9m��= �������{�uJ�i.����e�03���)نP�� �R��|��8�H���	�iy�{�O<��0T���r�:+>��g�9��~VO�#���j2t�3�2Y�����@��Ѝ�`,Q(��d3J�v�!�L�RmTl,�bݕ�N������w��5�K��ẒR���/�إ�G�h��q�S*�H�����'X#���U>��e��0�#�"�E���}"j�G�ǅ"&���=��{�\d��l{��tZr�i�N�c�����9R(�F��m@
�L��8%j]�6RT�����|�<�莰�'��sD��\�*���{�fۻ��4������];�p��Ή�KL����x������ќݗP��t	�s��X��T�Nƭ#�hsO�^2zQ��rBf���g�6G�F��|
Lf�_����|h��ۼً��"�<������>�F�ai�|޳���i؅��8!4�2�Y�(;��y9�����ĬV���c[gC�O��uF��xG��A[�`��{|zo�L�,��h(�?�a������C��Q(\�zn_�k_؅����50�h�m�
�:F&��5_V1U����V� ���g:[�v�"�����FiYR+�{�J�~��j*a{�i���\��@X<��|̲���l��k��d�������f3P��.����%�5T���#�Ͱx�����1~�5��X��{e�_�����~Y���7�u�l� S�f�ف��8�n�CC��3��Q3�AS��5���X<�G�(5����2�]1��r �X�A?s��/���!�(O����7���]/ =�Ȩ3 �g@���&Ê/�P.�@����L'ܟq���9ձBu;�K"�����w���^�s�<U)��z�l�r��R���[������O��#�{�]�&�^V�Ǆ�����/z.��������.�I��=�+���R�+\oc�O|�3䏝�������_��Q��u{h�J`�{U�����x��rv� �տ��2?����M܋�0Z���u�y�9�����ٝ�48w-1��P!�M�?>�?�h*QsW�X.����x׳zm�`f�
g��xc]w�W��;4��uF��P��l���F���H�;0�u�R���K�*Z�8�P_�2p7����?z!k��a/��|����/�*���I[1��x�e�l&������Φ���|�<ͺ��B��5��Ƴ�E��������m$�ۗ��Q�����G�$�d���r�� ��S����נ�,8���^�IAe�eA%�Pn��maJ�<�Ƥ!��>��Jx9�ķO�L,mX�h��q����wX���=G��T�&*.h�[g���r%vR�pK���K�N^a@L��ݹx%qa���Ǧ��^�^�7rD�/ôgy����Y��NZE���I| k3C���z$:w�b�9B�-�'��l��?��d������7��~g���|i1��T�ҵA���{!o�Ǽ3���m9��Åwm����^��*��'"a���px��k���7_�-�3��a��ƫë��)��.M<�7�z6}�11����Dp[��W��aM�#�+�J�NH@N�%�&�
)=�/�Bܯ��.�r8����;�J�/�9�c����I�⿊[������[|���Y�S�<����J������A4���k=ü�O����jG�s�y�N����>��'��#PrQ��l"�pHd�2^���2T�9���{.�0��K�X��b���,^�����6�J?ieU�U�+��)�� �v_k
Ѹ���T�*��jn��C�M��g��wT�[1�IƄ�PЇYh�tMR�Wz����n�~]��,�������$aK/9�Qfsh�P�$'5�Zjs���I�����l
��<K=j�"�I��j��^4�^N�'�IK�fͥ�m^���lQ8~�]����K3�<ӧ��/Z���ܲ��0��c��
�	:�ZW�M���{�$���zmcf[|����Gr$��<)����Orz�9�|��vwَ��stZ�~E��wt �0�!%���hAi�^a���4b��O�h����m����4n�hY��W��&Oپ)T*����kX��[?d�S�����J������UdDٹ���p_�"��[�W�1�+��%��-	.*�ώ����A���0�P���n��D߫������Z�#�����GF�7<Ț�l9�'pP�t%ɜ�7��lə�����V��A�F4U#i�6`, ����]!��g�rw�B�&��^#ZGL����j�_���ׯ�f�/���f΄?�9�<>��0�5�P�ey�)"���#��#�#�m��_{����4�@��љ�Waˊ�d�Ee�pgA׸-��]�2�����N�!�7ލ7᜔�Z=�7	�nM]ITӴ,*'Be��%*���<zY��YH���_��d�P�JM,7��30"�"���"�Zq�ߠ���1XP6�_=q�zҷP`j�M���c���(��r��ğ��ii.�U���_�0�����%{�c�j������"YgA�渦�l�=���x*!6��6��1��þJ��&��!���ٰ�{4�/�������N|���$�xu.�k㛈1�Ä�5i��R����~�<^^�Ug����H�\c����9��i�U�Ec4n���i��
�41��� ����!����TY��B�׳����K����)��!��w��T�5.�)$��d����1�S6q�7Ux?�m�<]��?��,�plp�j����5����%�.ׯkKhcT�s]�	Ǉ�R�NfJ���( �6�G��5�G��U���E��ض-WQ��mꆣ�%|�H�����?�X�����#U������A���-*(�56DN�.�H�7M'����'����x ��W�C���ׯ����D��
�$���S��`I�f@=leW��7l��0�j\�|c��s�_i\�~E��M����OL��������� �©�}ʞ��H�?��u.İNP���M�n�R_�r~�7|�zŉ SxE?�蔥T�t�eZ�y$W�����>G$�J"[�(Bx'>V3JR.�C]j�;v��&����NzpJ�4H+���<n����A�Vh��4R�\�'��^o$ ��gr�ޛZ?� �[��$�l�@�)��/���s9U�$���w�뾆�[#
*�.�z���d��t�4������*�g�@$gnῒ_�g[����P�\F�f�'�fD�`J����uM��	��v��1�;<�nb�Ƈyd6o/�+Ҩ�7��.�c^.ڰ��1�h�M�py�� ��4LNk5�a��[$ܦ��P�o�a�>���Y�+���L �����&����|�3�Ug����Mp�D�Z��N�l�e��V�>��\�W\�����a����9)6�RXDy�ti{����� ���X���L8·1��~4~�:�����Ƿ����A[c�!�]A^��5y^�����f2��c8fŴ7Fy�ba�N�=��	�j�#����[�����{�T،t��32?;n�Z+�r���Z��%�A�!W� I�}�W�+9kg{�^��T����o,
K�xH�ӞaupI�cE��xS�q�mU��y��F��/	u����5�rM��5���A?/���֣8>�eʑ�P]�Z��%��#����Jw!ĸu�����5�����jROƪ��]���	�\&~ GZ����[B%A��g��a�H�J!�������U K�������E3��M��@4�����v>�K��ohÜĺ`��j�'��c�B�E�w5�1��	�7����n�i�a#v�/䰺�݀��W�a\�N=��.`�V�U�LJ�E�ͥ���m%[��g ��xU�=�U.�ʟ�?�݂�w�e��I�Y��� �`�t�9$�A�¹l���PsP:�+����'�Z��5�t�Y?7g��d�|��g&ǯ���� �?��%�=N�bC8�}H�Y�{p����$`��#I8�	��0	'����{1	����l a��iL�,���4 a���O���}�w:��1	�tW;`���>h���i�.*���o�e/MK8-"�4
@���=|����o�g��M�UAEs���tq��g�Z�
����x�ʅp|K\�L�»���&������R���Xp�f���,|���Y��h��<������x:�~�]a���#�V�� �����S�flϿ�f����&̥���Գ-F��b	�?3�����(�%㔰�}�U�<�n��G2e�~�ٵ�εm�!(x�һ�N��$,o,J�}S��=���S���|�����y�F��RCa��X�14r�f���5��*h�-���8��� �з��a���:��/<���?��OK�OS��$��Z{+A���7��(ȯ����v� �}�!;���ˢdP}��%�|�4hY�b�Q�O���)��2%غ��%c#Z!2b?����:�뚽�Q<_]�A+�G6.윶'z���t���ސ0�Ϭ�4s]�"p�t^�w��=����١�|�c{�[�omڒ���ၡI�2���'�ٍ_�H��G����ҝ���_P
Rӷ�sD^4���}dl�l�#�����8I���Q�矐�t�}��<��+�S�?w��B}P��w�d�x_sP>�>o��9�qכ��Π�XJ7X>��>]}�O�N[_q�x;�uG/�Z�k�d��x����M)i{n��wm.\NU�S�����(��)�(a�?.��l�z�o�ɾ99��<p�իz�P��P�z��Ñ�}�P��4fdLqjzB�̠k|��H�SjwQ�t1v)��1Fk�L���?|z�5�j�aC��+��
X�l6<y���C�K�\���;�G�B���캿@��um�\p�{fS�:Z-%W't�/�����S�"UI��$,�F��N�l[I���![Q���Q���Kn������Q��Ypx�F#Рʹ�!�����<r}u:�_��&�/?P@��rgc/"��������0VSK ���<��z�F�/��c��B͵����O�A�:��9 n�����b���s	��va�~h #���m��3���8��&6f�\�I��M���Io���v|��ኊ��q�v�M��� ���L�� �x��~	�c�n����П�#m�͐%����{�c,R7N��{`��p�:)1�d�v���,mp߁'��	�;� HbE">I2��`{:N������4��l�ף��-!:Q�쳓����T��2�5k8u�����j	�3��7t]&�Ґ��B�o[X����xqU�!�3��M�|��OXd)�~E{c�s���e����Y@��-� 
>�!�Ĕ�oJ別^i3j&��x�"(d'`\(�R��}��l`��7�x�? @���<��4B��<�j1
.��!�Lt�y<?;�%����W�zr��e��5�w��W�~�p6�IGR]�.q���*Չ�%��Fy#௒$�Ulۈj��7�����?��ULka)$�VB߫�?�=$�JN�c�803t>%�7���L|��i�I�͡� ����d�,�o@}8�A��� �u��.�Ô�5�i�5\_���_䡊!_�q��| �ngL���	ݾ���͠x�%���6}�f�m���G �����Ed��B�_�m4�Y�L`�{������A�HmȌ������Kg��1�2�����,��;����`C�c(>��
f�C�t��-�F��Sא[`[T�
����� ik�PT��F���̣���s�b+qf��'�������|Cv��M"�y!8d-�����#�gC�U������_ �}u-@�%5�A�����I/Ĕ�C�|9��Sߝ�c"~��qo%[��a|���Q4�o��F�+ޜvZ@���:�WVa����6�GU�l���.ᵱ1���,,/�S���?j����	�b��Z�!�T��e~��0��R	�GwNb'��r���*�I�0��M5���VQIik]��-D���p��ڎ	�!Im�~��ʝ�&��Hu.��ؘC�$j9
�2U\)�*95}���&��o$��{+Y�W�9�,�%2�`r�L㚛 $U�
p�"R>}��Q�(�ߋ&�k�����Æ�C�K������>�D��*dX�Z��s�O�q�����;���rJ��m�p]{�$���΃"a�*�z�cg��D��!��:H���t�P��M5%�D ��L
^�#\e��ѽ�R3x.LGGA���U�p�Y�[+����K����!�Ά
	H�qc58@H�sLk�h�w�,t7㾟T-k��w������%$�ZwA�/ӗNK�{�i��щÌ��$i��>���)��w�:��=oSs{,�£_)�/���Γ��*��k! �E�T� 6�����T�&r�`I���˛�# ��ըI�"�~Qw�,|���t�C
@_C��:��|(��V�`�8�f�`O��`�?�G@/�0ƥآ�X}�|F?vj=����^�t�����~xv��j��1P1"�ӱs(�C[��W��m�_�QNH>w!Gp5ӵ$D�/bB��?�!�|n�T��RF�d�+��7(v�w�6YX����{>0����7:����c=hTP8�^����F��N�m�H$�D4���܇�2���66�߯�+o�����͋�')�Je"@v�L4��p>�����:T�6s��.]=HV;ޕ��*	6��I�c'�e�$�8N&~�A'�=��u3b,D��pb�dY��O(�J��"'¥б��wv�����/��!�1!����K���`�*������BC�;;;��8�02���L��B���1Q��@.'��MMVL�i�*eHs�;e�z�oX(���w�-)V��`�oÝSq�S�^��:�p�X��Ռ��-'�e�溛��l�r�x|��=��p���G��{ͭ��I��|lCCG�0 h%�>8�K��e�]\�͏���ү([�*������7�e�w�Ĥ�öJO���%���d�*2H�Ȃ  5�Q��Фu�5��2)��c��К����Wf�1*����nA�YapJ��ئ���ɽ����&j�ͽ&dЩ��p��I;��I\VU�3r�a��J�&�3�I������w����Ӟ��Ƀ�4�E��yap�L9�m�;��A[���$�8V��˛�*��5�!,�)�X��&�VP�g��>�ӗhܛI{��;a�rP��� ���2�2�EnK��O
����/���x�d	�#P�S~ą���k�D���?���do*�|Sƛ��'�	���
iw�u&I��
�ѧ��*5��M�����a�ȷWVvkSa�"�O������2J�gk����B����˯�.�oe�h��[}��٧�.��<������ kD~)��
�����g�`�5	Xtrg��7��������?�*���6�����ԍ���>�VUA��"���K�R��r�Ip�ߛ���mѶ
�8��bqt��D3� 	���4Ữ�-�
�z�Y�%^#�v�9�sj�f���%km�P1Sˢ2K

�N�0�"�9씷.Gc�P\�-Ѹ�d��"��i͞=�i�d`~Ӂ!���e!�٤{��aw�2��� ��N��=�O
A�1h;��#LS�����\p������(ԝ���g�M�v��z���N%	�뢤 ��~"���:\�&��ը�5I�1DX��q/��%�����K0��|/hmb�~6W͹{��{���p�,�H���q�ٕR�w�K�OA�xB%g����R�>M��(pȃ�R�B�K)�g�����{���'M�ei�M�A/B�f<J�<J��m�]>b#pZ�!#����ܷ�%��"���@�4����U9����0���P^		��s|��^\���������ߥn��F���b,���� ����d+�{o��"Xl�BoQ���h@ZP����� �pff|���=�ع��5k�S�3��3�'4m�If߹�}<@"�~>ww�00�1�rO���S��>=^��9���D ������
d����Ԫ�C���3w~����|e�*r�1���9``x��mFg�\�iA�n��)��&�\�ڟ}�-���v�M�N���b�Ц�{��-Ӡ���-I]�(���y�o�1Cܵ�qy:uǤS9Jr�!��C*ŧ��.dȚ�����a_3����2�� ]��*�����h3�lS�`�`�Q��sNLB��$��z#�~�s6q�a+Z����� $ei����*3hGV	B9RNHJ�Cw8���^Ȝ�� �w�u@��j��&M��ѳ���pG"�����ϥ͚�Y4:��p�o�J�E:�rY�4<�$��ݹy?� 2�*2i�[�e�$q��J�$w��[�\dͅ2��f|%�)���H|�,��추��}�9��ս�NJy	�=��:V�9@�&chϕ�EL-Rb ��Ms$B�˙?��P&}��P|-�j� @v� �H��M��7�d!
x�Y�S&L2)�I�r���hpb���{a�I��|��Y�k�^��
��ۻ�%\��j�<�!x�ߩ��'�[P�?ޢ���9����Ѱԁ�{�4jPٿH�.�S��I�%��]t�"`�i��;�6�>��g �[���ʢ|G�fAp��ئ�u�tA�2I�:�PJ���3�,��͆��1���#0f���~��*�X��G �v��c�z(<�C9�&O`	�?ׂ��=d�ٺ����F����r(h{[��Hԃ �zx;\��)ʺ��o��n�M�k:?@�!�c%dո�
&��M��6Gʹ^�Ƕ�c�m�?�i݄&<�N��'R�_k�_�@�:~�����QA��{BeF�t�e|��̤}.m���5����ʡ���c�n��T��^�?��ѐ3���"6��7i���̃��5�?U�C3h�-5ݗs;����̆D-�r��ѭ�S�_$�aTpD�c�63��N	���WZb�zG�!�r�#����.�#�{+'�&���Ğ��A���׼9��G���'ό���T�Hh�Y�U���n����Bv�ԔJ�r�����Ԍ;g�>��3���?��jI����Aj�b�T)���,{�fr�?U�Q�0�*_i���9}?S�[��n�3�evU5�29�� {M�qH�l��F�ѩ��pn���n�=pJ�#��2���/{�ހ�ɟ�-��&�X�@�(;�C��D�&�Ѻ�nkT|����Gݧ���ly ���՛��U�
ۇ�l=
S�S�,lqm���wA�Tp��i����j���'��rP4� 9s��M�� �k|�U#J���]BB:��$��,Z�?�]r�E�JI���Ͳ1���&��>�����B�D�Af�G$ M@"ܴ��&l�b����=h3:����p�w�B����x�x��92@��� ��9~�i ��T�\E�l©��[��kιr�T����V������ߎ�;mm�eY �z����`�_��N��9,<��lتt��1�zjzň�|(��\���.;�(�*���4�d)��g��z����o�f��u8�J@(V��������{`XA��"�gz��B�&p��:�F���V�[߉e�:=�����%OO���3�>�at�ڳ���>��]Pꘈ���,E�1}�P~��5��SK
�}�p�8���v�n-􀱻�7!=V��ͶJ���VZs�6�F�kF��'J��)�@7�� ����ݦsy��ׂ3}{����n�9�������U�vg7�k�< �j���Í-�`\RӀ��;��a�u^')��NB$"�K���*]B� g��4Gd(��d�������M�4��[m�e����+4�7�-��L5)�:-O웂����p�''Ѐ�C$�M�����p'�0����r�?޷�����Z�AR�� �
H$��!���̜n�_uғ
�|�S�zO���1����n���ڂhԡF�^t���Ϧ����Up�t��g&X�� K(��zE)� ��alV�I����d�\��j��$��V� Z؎󎎏�?�x�05���fWj�#����O�_Mڋ�� Q��R��~3y[)���ځ�յ��@���ho����_<r����Dp�MS�oɝ51��xÖ�:�J�Ts�����`/���t�Ml����p������
��{��2e��R� 
�~E8�ƅ��i�v2��kh�Y�`�'��#�z]"`��$�N�n��u�M0���5J>$���� 9���0.��P%����K��Y��T5�g� x����"V��)������6m��n�X�z�\�@
%dWzŗK�m���L�k�T<�@����5U�z��:�*��+��c�Sf���k�������PdM����(�cǇ:Du�x�_ �_<"�<A��^���m��"7D�t�.��9ǭ� ��e�fQ[�^]Ȼ߫*r>U��%�d�iԣ�?P]y�Al�5����(����-#����}&t1 `/U<�1���C�|�qK�b��VX%�U��5��ѕ6ˢh3Rf�
��2��z)�zD˄�����P�<x��E2D��f��7FZ�c�Љ�#T�J��vi��f���������	���y�=��Qv�@r #�qFqS4����͜�4��$w ׸|��N��h75H���:�GI�8[Tv��p�g
�_�Ƹ�Tp x	�c��h�y�dǥ�*��L7��µ��=Оg�C[2[�~�����7`) ��Wp3�c=ɕ)��%��z�+ '�x�����8���D�.5܀�W�y�6��W����֔��O���S����R_�Kؙn�ưJ��%Ĝ�20�d���H�b8}�%gu��5b�"PD��'���O桡������w�*�qʶ?ÚV�RX��H�E��kof'�SR���<ԥ�<�[ y��&�W̝��>ʥ9]6�~�Nٞ�r?��WJ����aZcO�ng.M�F��֤�J2�RM�����qCV��F���c?��WOq�c�Z�e��<��s��]�3��ܮ�:�+Uc��1EӀ::�?&z����b!M�Y�C�$z{����̨wΙ�WZ��qu(�������l�5�]���3�c<<{��Hcy2�����sg8�~&AKъC��C?��E���ࡖ���ZL �D�R�F����C.wzY\T=雵�O�l�!u�
��e�~��伳�� {Ƿ@�O�G&ږ�V1:qfʵ�D�Oq����g��^�h�̭��f����+[�f��X�� �C��n*��ѝ�-�6�U�%��!E$g[ߧ��p�`�SC-�~�-���ț_X/_�tx��D�x��b���z�´_���3�I";q�q����R�_�tpeggP@;H����g�֫ �N�4�������(�t�D��X=����zH-��Ъ�&��~Ѓ�����2����s������1H^05rͻ��0�^
}��.�~ƌ�%v�V���EhsK߳��s�xӕ!K�I�Piϱ���E?E�AGX�#W�Ҳ������!Ẹyv��UX��'�#I�qe�ރ ��J#�$˽;�4n=B�M�f�W�xޱ��S���.���� IM󰤣Ϋޕ�wLf��+����� uȕ���r�d֭ȟ����^ P\�#���e)�mR�AySa�7t�H�A�L�-�Xي��bE��x�  �	e��=f�z R���	ߋ}��#�$�[ ݴ}�b��1�|t'$�m�W}c�uXl���>������i��j�[?�Z�X���X�������&Lac�g��Ķ��u�a���|<5m[㍼x���E�afoȱYw٠V;a� �?�]�^�8J!I�pTpa <o�+� m��do��:�P���Rt� v�E<E;q���Qх~& ��e��1�DH�y���X�!#�{+izA�u{��mk�c��#T��R&���$Y'���P�J4�k�rU����E�Z� �x+�=��5%AW!�_�q�4t�r=$�Y���t��5�(�y(n}	꭭�SfZ��6�ʚNhH��`�V^��}����`@��	<����> W?�:����J��{Yotjs����b68:��p�R��+鼖���FD�z�:�?�J�>�q`P��m�0��-ߋ�~�X��w�$^�L������$wk���$�T��y�7n�ܠ��g�Fj��s�T��`�� (U���_��4;����#3�,���Q�u	���q��3��sO~'�u؟���)�'�i-�N��a�� '�ޅAW��@ilb�>��8ٵ�T˱��t.��<����]�m�0��>�I�M|��W�5�S@t F�R�)
���Vg��y1�:enq��Q.[��Y�P0ǟ�AY�6U�i�@�J����9�
� @<�ޥm)����A$��^��5�G�K犯w�f��ʐ�@�&�H`�-�{R��ޞt�,0Y�� W �Lo�C�?�Am�i������l��+�y���JP��nj,4xZ���q\G�^j4!���H� �73�6P�UO�����
U�>@!ͱWa �JL@���q+�_6d|�x�g`!���c,#b��0F���^�d5�p��l`��̓�0��\W`1aWQi�\-E�Xc�ҟ�KΦ6��E��
��H�#nNR6	`���#4o�}�(�N��|'��ٶ�d-:B}54~\�Pn�g�V��\-	?u��˭���J��=�-������f��U�-:4�lx)$WN�&�����Rƴ^d�6�6h1�/0�p�#�r@ImB�-ԩlmD�lI�����N�����۴���`ľ�F�bW (GC�B+y&"r�����-hN�=�� ����/�u�5�2{�3n>�r��rQf�W��&���
.4Y5n/��_|��&�^�
�N�K`�ȱ��_�]�N��?�
B��s��=ɭV���� ��(�f^p2���}ǍS�
��T��ؔ�<�kX�5�;L����I�_^�.���y�ܑd~�Pc��y�11k7��7�:R��A�B�ˮ O�ݙ41���#��p.m3Y�P�R:W�[&S�>>�jS0 ��h�}�݁{~/k�%�h@�S��r�B,)�;j�ښH�� �_�N{�4�S#�R!��F�}��d�P�������vД��2�Ew滲-��.l��9���9p
jЂw>�8�E[��r�5�K��Vg�vOy�v6�J�,���X�+��:�V�����ͧB�(�A=�ߊ<�V�h{}�J�����zw&�Ԩ�-R��IS��Ky#��@m���M����C.�מ8���b8�V%� .0��]�%*4ot�K��N���p��Y�E��z��EL��yG'�ۣs����J	�͖��K�͚	�9�()����f���
����7�����潣n*�sx^�D����S�q�_���|p����������C���b�c����Zh����kZ�/������;j`�5�Τ���/́�:'���\�T�naCݨ������]���݀��Ш� ��4m!��)��J�?�q��1Xt���۝�7|�R)+N��|��.k��w���uahk}�8 ��o��H�5u  �s%���d�n��3��qe`��s�;����	g��{�'��!p��f�|2���,�F�}��ӄ"?�b/��9��u�?��xF�x|�۩�\����k]Ŕ��#�'/.tJ9���o�w�m_��:+*�Z�ڨj��w3nJ�
�����ް��>s�ӹi�Qs]#t>�֡h�V~V�Ύ����J�C3���,�P�5Vc��ۻ�B�+;�K�nwh�Z MK�+a9�ղ�Tܘ��{�~�����ߧ�T�;���-�m���&1R 1�Еo*4^�¼;!���x���-�>[K�B�#���L֢���[uO�3�?��~O+�\R��,&4�� ��ky���t�=��h}��}晊�ɞ�R�*��RE]�2�:�x���4�
ͭ�k�x����v3\����U�+�GTH��_VO%�~�-
ֱL/^^1{�d^���T%�˥�|��
�ZYh�\�<?�1^��c�E�D�C�Y�P�5��/Ȱ��(�}��TSJ�%P�=s�Ȭ�>C?���_(9D��>ܩ��#��a�Xލ-#��:��d���F���E�M�(.UѺ2�#�`�R{�t���u%����j�]	LS�B]z���-�Mp���~����k i�'�(�>�ixW��%�y߸Ew��;��X�߫������3��"a_����d �r��!��?i"�r���PA˭�$�X��4Q/4|a�n>�p�O��z( f|M	��#+z������X���z� �u��8`�!z��|ʞ:6��K��l^X���Xh�n�gi�_��I�GR�0��{u�!uCϱN���tV	Z/��-��.�o`�B�E����U���ec1r�ҞW�?_E�>7��� ��F�l�vF�=Վ�F���9�B�����	6���}fĞ�%L�򴒆�jϑP�ę���ޏ����� ����Xd�rV�404t)O��dӜ�è{��%�ʍ'_X���t����؉2[v7�o�U�F�aX/>��:n��:�2�y�9�.���5�;�<5o*�ӕ"��S�)��Дq͙D�tw��R(GS�����$��8%*�!����^G�ɾ�
��6����9�6��{�5��`��w��T�4$Ò�9��_$\�i63+�V���A�v�-K�>o�������T�\ڻI�@o��&�B�gW��V���+3�a�W�l�WQ�/�.�ڦj��X�)�%��6�����ܖ�ә�m+ʾ����xXQʣh,掊_`�KI�c��̱�Z3�~v}ʴ��O�����=�Ŭ�[ؑ���譄֌���^���SZ�������<+���	����og�����1����Jy/�^6�R�o�j���`��n�s;���{z[(ә,wzZ,G�c�(�=�YJ
�k��zph���T������N�ZD�m�\�ӱ`u�b',�����K��%�$�,F�w/𸴵�-�f>���WS��>6`+Z#\3����J��I����am7��K⼣��^�k)�pF���G��`t%���d*z՗W�!(�,��N-g�+��e�L�ٜB��9ᛸL�Vie��-�&z�����f��ѓ ��LU�N��bh�T�Y�k핲���+C�U��0?�'�!r<pW�c"P
-��Ni��Ḝ�����%`ŝzt%���H��2nhz���d��Ħ��QИbpSG����3�q��v՞�����\��.�T0+GKcb&��pw�S�N:U6���x��2V�0�^�A��h�Y(	|G�$& ��5�`ҦSH�	�#�	1��E�)�L ���X�E�������>s%��h�<,�Q�������V�>*�y[�ל��&��~4�ՠ����g�q���ϕ(o5$�Rb`�׃XЖ�4<�0�ٰ���4��@�T�I��Ř�eq�>g͝_�:?��k�9|�.-m�9����.�1�R��í\ѽD��z�L0G2z[шo1}IA�����,O�T �*�}RñFQ�M�������F�Wriʩ��ǝ��݈�P��̝�LA@k�SE��i�G{�aakj<�ê�h���S���`���)VS3}�R󰾺�1^���� '��j��7�bMx$
���c����oڰ�B[�U��Y�~�$TO���:
=��Ҝb�'�oT9g�g�Z��GD�q�7"�I%�Y���l9H$���+�]+B鲥�gjx���6ԙ�*�.����|r>�(�V'f��T��R�ĺi-d�,p��feP�wI��l�"��@��yV�m�yS�Ȱ�s?PRHܛ��kg]o� VIe�jl�)1�J]6}V|)��,<DŃ�&�h4�C�:�h
GK �:@g	<Iў���F��xj<�3���K#�7)Ӵ�	Y��O/<"�x�am�v��e��Q,�Xp���S�.�9�������%Z�Q��"B�r��sx���*�t�!�:%�)Psgx��A_�����^n������J0����7�W̣,B�W����̝[�/���/P<�+�	H��������u^�y��Jg�Ȋ�;}q%߫D�܁V(�TN$��z�\�{Lx.98���]�=|����C���2"��$�"TiI��Gj3]R����H��:)����%O���u����ѝ)�f���#Ո���\�p6r�2<!
i�d�������i�@z!����bzw��y���X�oXt�lCE�.C�Ԙ�Ĵ�t�e�w��ѝ����PTL�I�[Q��ьt 1�g�yF���ˉ�h��>/�N�2�*k��C*��Z+���C�OOȫP_m�?��B�rW�(Ժ^ײz���F�����r:�*��]��ϩ�	�'`�_������[]f�E��w��vv�U�R#ǻ,kiǰuM�
�an�D�+F�S��<)�]6�����#e{-D!5�i��Z�E���b(ӽN�����.�_�\�,w��Vr�o�� Żb�[��3m��H���`��Z������u:1?-���%�������qF;�nM��yg��2�c܁��m:	�d��__�P�^m2��4�L�2����x�]�^���+�v��^�� �@$�k��2��@U$o`��˘�	K��O�֐�s�Q�W�Va�.x��<}^6���@jG�x�N��x����A'��KM��"�VF!�e��|���f\u��.��(�K^6.��c��x�J=).6�1
�x�z��,p>�<m4�dt��9��a�&"�n�od`99*�o�ݏ�Y��[<xhN�������9<6m���)�my�NH� )���c�y���Tnus��J$r��B��3��~T����I,0M
6pwM�`�˞AM��欥��N��^�s!�)��C��pZ!ڕ��1	�M�7@9�3��k�M�Ba�+e��i��9�-&���"(�=��˨6�N�lMQT�cs���#�iXk��QQ�8I_��d9w�80��?������Y˧�3�>�3,��4^Ԡ'r��Z�WFzr��|���q�F�O��Ou��n��1Za��N����\����cf���y�;|��d����v"B�~��ؘ�>�<Hg5��ի 5x���1:.�x�S�����l�a[��|S��/��[��hH�!X�
 7����A��Ӹ�.9>i�],ם�?m:�56�V�jaA�<��n#��S&(aS����}2$����Gw�1�{��^"�Vi�!�%��������H�A�Q6(u5��>���9B�}���:��l��̼�fyrD+}�ۑ���)ݚ_Y(-R��i^��ǹJ7��h���%�H�L�?��,=��|�.��ȱ�ez�$û�T�B0M�g�V}Vh%� !��qf��%jwǥ�r�[9���
��L*�Ŵ��������]K+l4/�D��_���dN��=��Rc�\����xV��Z�Ra��ߜ�.b�+��t�����[ݚ�^"�Q�Bކ���g�e�>��[��d4]Dk�)����X8��xv��o}`��^pϹgt��G�e�!ә��NgG؊��eI�ʝ$Z�qZ���k�7$kh;��(��m`	��\���8��H7��6d��	���rw�\���/��~�����6��>��9s���1pB��j�r3BW�;�bò���^���5��9�.�3U��!�����x�|���^���?�j�4*�I�8>�k��摚F֭c�����F���-*;�����j�s����7N�	�	�@,�M��Ŝ'C��η-F {|��иEk�I��Y\~Br�l,@~e?u�]�V��ٝ��3߹���Ic�kF�FD�z×�|���O[K��Q�X���t��s���[���1տ]�N�ki(�n�ւ��o����
��Ϝb�E)Ե�i&8�|�����}יͯ�����~4W���q�eow�憌z�ޢK�3_��񧨭R��<��l��V�!#���Q���R�U_�D�����5�0&;��=�<kG������l�e���p��΁F���<E�;~�SE�i���S�z�=�f����4?H(\���\�_�o����*��좬xڞJ��������{OH���Ɉ��	�e��|��	�͜5yZ��7m�?����'�E;��d�>AR�T�uqZ%-o�����M��/>qOa��%���V��W^�ҍx�k�(J��y�qˌ$#��k��R�L1���&���,�e�ٯG��T�4^}A�f:2��
h۪0��]3��m�c�����[���a��dT�Z��y�������^5�EUfr����'�J>���	�T�ڞ7F�ǆ#]ɲ;UB�F<����b����Z�nF�巐,����F|��?�����__��aҁ�R};Ƣn軆��t1��fDl*}����֟w���)Y�����{6:�;�Ȑ���w�1����c�z�?�_d9�d_�5�H���Ύ�N!������*M/d�LA�T��<JuxF�P�r�PQ��/'z��>�m.x��4���rՁ����[�eR6w��ʛMډ��;���w�7<��S�<�\\zJ�&{ǡO�������/�z} I����}��C�zшL��5+���}�<�F��m���P,l[�{헑�O�0���.�9�$�Sp��=�k?��Yoŝ �� EÅ��S��X�̀���͆'�6���ƌ�]�������Z7�����Y��ܦq��_�}�j�s��7��3����8�>���~�h��	=�,�CcU�}�O���+#Vp��8ա�MN�AW��k`׸��{*vXؠ�Zpv*Oi�߉�O)݈����@};'-z6<d�ڴ���
�o���r���ڭn������i�j��\�/���=׌�W[.A�d^(�E������[����ڣT���~�y���T0�O gI�h��-�KN?a�	�|A�Ghwk��M���N�7���l�P?P_�����#z�\?�Zf�NR�3���{����;hh�!�3����� {�Ks4��[X;������V����<y�$�w=u:L���̇�������A����~J�ޙ��糎�c_�,wj-+ls�c�=`��L�oKsi��"�x�ݻ�v�@d���F�3sv�B���S9J|Ď�E�5���,<!pE�\H�U1̥=����2��1��ma��Z����~¥!*�Jb�2�:�e����4�����a'�N��8et�K��K�p4�c�@Z�l�����~�*����3�tF:����"Q�_����}'�������~:9�P�=��D����d�O�M��C֥�vZ,�\���|r��Mn�ڙ�!	�z��󒇁r92Ux�1n�m�8_t������ʹ�@	��d�'�;P���2/r
�/�EE��~X�Y���m�8�g�`X7�c|���_ڤ֩���$�H�aа{j�����F�4_�NG
���]g��e�wq��8^�C�]���4��i:T05)U��U��O��=��H%4��t�!����S�Cή�sU_�܈� �a�w�kc5OE�ʹ�<�%���
�����}�z���z/(u�Q�گ��^�חp�ԏ-M�p~������J���x�����]��w�'+%�U�0�?�jU3s���CQ�h�g�&��̎L�J�bS����@Ce����Ye�E��F��G��U����1L�Ѷi@�^��p��������o��3�h 8�zȓ��oވgtT+#���v��@����+��A��i��3_�@�Q(�v����Ѫ1�����W\:��Q�Uo�9��v�W�U����K��rVł���t�tW;�՞�ʝD4ML�A9��J��s)��%w�Â~p�̝�3}Y��ހ�EY����wG��~���,���3��	��v��i�D��GN��B��!��U>��od��[���	�����m���6��~����h����Te5.j�9��XP���G��U���Р.�6����5p">�� a|��-F�1���s*Ӡ�YA��АW{U(��|i���'����?�'u*�
boaI������?�/A���{q�Q� 6��*uҿ���J0���4�2�riSşm�Mʾ�?tNuL��E1x>y�/��X�3�P�|>��?��K<̸>�m�r��a�<O?���$��M�D���l%���#�[F�)k�2g&���<�7:�p��u�Va<��� �	����&�tb��m
���m6���Óuv��Jq��� ��y��c
������!B��>@��I�H�ܖ��b<EmG]�i���^`�#��Ǐ���|3�DU�G�Te��s{�g������q�O�D�����]rmr��Hㆿ[T�ȁW�cQx4�;<����&�Ᲊ�!.��O{�\����ʸ�o}R��B������g0�;?�pR��K���aD����	*ǣF�l�E�e�������#�Ӫr���dP��e���ϱ�@��z��z�K����W2u�}`{�F£�6T�ڈ�ZU��GlR���̊�0���y��XH?��m*|��x�^�7�D�_�#�/���Ar��A�_���I�k�W����S��N	�[on�����?�ϒ�c��n(U_3�3r��M��̽�S�{jw��Q,�<9K3�M��ڞ�]����F�m�ork�x����{ӔX8	Eڤ��D�����z��0MJ�~����}���̽�U拆����S���N���V����{�,�%��{��G��'����Ny3$����R?��������a����X~GP��;R��s���J���!��kg�&5ǡw�<�`���o�v�'s���5���k�P�~� �;םS�>�0\�����DL��Up�/��Q��=����%���D����������˚���}.;��w�\�	ioЭ:��v�+�"1��`�\+;��|��m�D�f�gѷ'	ܢ���Z/�[ c�"t��c.��;���S�k��4<t�$y�1>G�%���Qr�{ȢylIz�-E�?G	���k���(g���Eh�TC��/GP�l�3��P{9��9������>�e��ƿ�:�����'����O�$چs#�ی})�%���Lf�$>���03<�v��mK��>��>GU�(��Ak�ڧ��O��X8�D��!m�l���1z��:�H9�-L����0x�w�o�qG$�*:�Z_�x�7�K�J���t/\��B���wi�&]�$����pu�
���s	DHY���R��d$�[F�j˛�0�x�F<���7W$�ä|�X0�͂m�ˏ��qG̻���iE8}�����`����9o�q��3_�|(U�*�օ�(3�Mn���"��g�V�֤A�$�ݨn�v�穅�9�Z��g|ޜ�x��Vy����l�����ُ�d^�e��F�/8��J�n���l���'�0�3uv܂�Rm1eLW���>SQZO�4(9�;�ֿM���M����'�d򟐩��7��_'���+��.S����9�x�����sQ�.e橿���d�yJwI>�pXs��PC�aǫ���2����E+����$��J��㳫����Wv�Xt$ݡ������Z׮y��5<R�x�ɟC�WW�ܐ�Zƨ)İ�(k�k	Lu���Fi����p��d��ɠ������M(��]�#r�~SM��	L��E�y���
ZKi�A��9~z�}��;D! ɛ�{�����ޕ��.U�2�ԯ0ye����8\�,l^8[���1�{��"��J�/9��"��"�\'�m��&1L��9�<��
(G�q\��`E���s���P�:T�zx�W�+¬~{`6�A��4؟���qM.��5o@/E7١j-�T;[�&�q�-�Ak�͟�C����Ó91�`���c}�FP�Z�^m���4�v����d�iQI}�z���ÿ��C�!�y_��/�V]�/�=nJ�n���)=�؂�R�^��W�x�F9z��s�l?`�U_Ӡ�|��?�U:D� ��@��{����%g!<Q�A�����j2aT�!Zf̑��y1��6��25I��B|M��4Xfb��M�9�h{}J��t
}>���1X�	E�!��Ft"��Wx=����I;�U��jy�h�.�|�
���;k�;��5R׬�����.���v���������_�$�~�yf�J�^�S���5�W��Nf�S��/_/.+cNMM�4�h�����q��"�������e�k�[@��MS�Tn��I�*)*�|��,~r��+���_��si)x�Z[[+q@�U�E����wFc�C͉ol�T���ȅ/%�(r���87.))i���쌳h�o/������C�e�3K��щaFy@X�֪q;���џ�F���ˆ+Gw>�������fgei��q蠩l�pΔH&r�������B������A�v��I�A_��,&+#�aw�hq�t�y�=�9B�؂���������N��N(�{�ʘ������v���%�;���эV�u��q�<�m��4���2`;�f�x�䅠�)�[�Ȓ�J��KtOq�f�N��?:.��K�!��U?U`u��E�p�s5��Gˇ�.Ec��Ԥ�O����4��)W��(�+`Z�����i��V�U�C��vx@k��b�M#I�{L����!�A��h�l��:ʣC��5��[�=X�)&ٯ��A���1<v�����+x���Ge,w~ �F��Sf>����"�o[���jB�z�|V�|�����wHC�?�-�	.���+�����e�HђKz��?����w��d�R��zG �#mk"�v��'͛�.\GPA���#�?��v���sL���� u��թc�@//�w�!�b�n�#S�����u*��'�|�X5��+Z��;�^-�h1S��%��B`�.B�!�{�Fd7l��=�S"!. 0�1��/	�0��&ɑ�䬓+�WN���'p��|-6�+mT��WA��[����و�Έ���q�O%)�$�ڑ*&0�/�F ��h� �rLN\���U1~;b�y+M���wD�T���i��y����u��WP |���� �R�I�Nj1"��ыk���X�:SGt��{a0ó������OLZ,�iz��D_�O��'52�l���td"
x���������~����)��@���(:��#�D���B�����3�t( fF' !"핂Ҫ스Up��:5( �� ���q�v�oc�Q7'q8�T]r��	/p,q�!9J��hը����3F�w iP���D2��F��x�<D�),i�,�����՚�͎Et�M�԰0.>t�`�u��O����0�����/tP�6�o����ԩT�N�����-�.��hB��kt�вګp�7FI��ź� �����~��u�h�<�34T�B�������:�>׼���UG'�3�- �Y�F�����?N?y�D�����b�j`�V[5梌��A�K����ccJN�O�݊��mO?k��Zs�i�g�M~��v�G���DA��(T!�N�#:K>��8(�鮁�lk6{r4���#�4�J�|�=?�Z%߾]�-cZĠ	hߑLEZ�h[�AI��T��0�Ù���NM8�N&��nу�O��2Euy����uT�J�i�Sj٠�s� ��J�㥞��	�Ng�/�}K�n��)�99�W{⟓�M��ݯDl� U{��&~���Z� ��(���ǜK��?���o�e3�=1�<&r��jaKgEÜ�.�a�o����Pz�|h4r꧀���0go*ʺl'�F �ڋ8"x���k�o��*���z��� �p�9]V�f.1Ul�Q���^X�h������U�2����
vS?��U��5Y��eu(=&�o��g����TGB�T��6�_�)*!��
� �sٔ���������'y*G��Y�A���P"�@,��/�yD����J����q�$��+c�+%E�ȱ�hgr�4$R~�KS�����*��� ���Eʕ>��H�Ne�f�g}����r�ؘ��ġ�{�b���a.�վbXH^ X��)�#.�kXnL��e)@�.Fr�,��+�JɎ퓉�eA TوJ���d��	]2.����(��c>� ��1�܄�7P /xY�IT�U��=O��L�\���}���O諾�XYpUޔ��j���W��w����.B 8gg�N?9V���G�1�W7�~đ�s��	�%���b�~���OG=����V���+�h���9�<�^l�V^��1Έ0UL�x���5f��������O����5������χy�HH���7�b�X5N��<�:�YYu��i�������Y��jsǓ���}�!Y�3�.l�@xSP�?���g����9�ޕpw �,�(�Tj�V�+DSk,-@��х����D�<ԕ�lI_�$���dBJ`+��a|T�v_���t	T�_�n9OQ�5��=t�<�,x\j}
i��\����4��F`Z�Ӛ��â����x��sT�p�*��	Siv���$�]�v�G����X�Gp��^�w� e�9��q����w���Gv�ǟ���qM��|P��RR4��pJ��	y4"��s�(�2���1��	�Ikh�(�A��s���>��FH�_�g��������ѷ_42I�Dw�H��x0m�9�kK_��4�\���!���Sx�s�]\�}@�4��7W������6�����D`1|�����Q8�%�>8F�)wcr�hk����:n��M�tI�	3M�3�t{')�t�z��V�	3�[VM��̴y���)8���#a�G�i�6r'�}1Z-YhIv�4�}��a������'ێ��O�<�G�f�b�c�
�K����k��<8�����~E�����'��Ø!'/�w�4kq�Q\K{�ر�W��i��/��(=$̍W�Y��נ���1�$���?�!`޽av��w_܉�զhF�1b���O)�E�P��<^�(��͎���*�x����7C!u�c�ku}�$��_�r����
�Q�-��������2�#fk~���z��g{����^�0[}<�� �_zu��n��9&�Y�q엤�#�/l�}�4��/�G&^ׁ�4���}��vb�z�X�߿�\�l�2]I�T$��C�O�O(�����-��ᖍ�����A�-���m��=�ֽ��E��!A�W{׏G�v���)�O�����~��l�u�_<'��8�յ(5i�ْ��^��.R�Get��^;a!��p/BBs�;�9���'�>ۃ�m@�i)NDY�QwEb]^�W}�ŝ���-L�G5a�[��gy�����}Gb5����'1�x!���C�$���c�4���M.(����u��#ǗIᴮ�k�����	ۣ��C=��'�T+$@�h��l�?���DS���G�`����_�,"_�$�jձ��8&��q�%�Q��Ɲ@�H٤����ax�ջἂA��Y\�$ZL&��)����` ��Y�ɍ�V��>���^��Ͼ�>(�4���3,�
7�<vp��0v�yp��(E#��]�lBu����3�h�#	'�r��m|�}LԹ��P�ҫ����u	������+3όc�{P�� �������/�Q�$U¥�/2���|nd{'��ـ��BM��`��oI/5���^��֓6�$T
�=�r@t�Zh��tM)K�{��]�*wo�#+�@/&��I�нNu�?"dw�UP-Xhf�������;X����Ŭ3�B���q`���	��)f[���҄R-�����2D�U�-y�7�z��<����IQ-�u�rY�������|M�E���A�D�0�&Н����p!2�M�W�2��km��Z ;XK����"HC���|�n��ˤ^n��Y�n��I�jڥ�au����I�&����B`����N2�vZ�����������(��L�J���Ȭ�Z�T��{��=��G�ӄ�Õ�~��e��[@�K�0-6AU�l8s�쑪�'���:������j֎{�Bڰu%�����"�w �P�[ʅ̨�`!b����ӿ�r<�G|�;>��z��'��$��ًT�#jT�·��S�1[��k���Lf�O���\m��ғ�;��|&��5�^���l?��mA��wd�V�"�K�"���'����BY�HF#���]QW��h��z�s�bq"�Gt��h��R��z��V��IoQ�!6����Z"��|�=��Bt�y���ҁ0���������#�/��R�(���7�/{��hn�+�
�k�zB0�Bh�;�=�\<� �Y�/����Z��LJ�ƨ:%~xv[힨��]���«��8x#l?��gߘ�0N�KMr���u��_������ZԴ}-���N40R�_�`��o"�� �Z��3B��Oj��M��:�.��(:�E��]���2�>,�^�ޏ��T ��ċ?��!��Ȏk��Bc�ф./�J���r;�Q����|Gd�)���)�-l��4��xf{�)G��;H�@�9�BS��QL��� _)�?�����t�i�e��q�4<Q�Hy����?`�<<��gUP(<�NY��F�_B����|�y�J-y3�q�W�"�O2Ǔe��z
wn�B�Tgc�e�q*���u&���7��!x��'"�c?�e����ۈ9܂-����6��u�^Q:�q]cl��+�B�.�f( �hW���_��ی���O��9Pe�[)���c
�}[/�Z��ӟD�B�p-�M}﬎@>�u��3��a�&�蝔�S��mxgn�y�m�%dE�7����-�ޯF����8�s��׏��o�K�V� gs�-w�p�'C�8?}�<��o��_ș���D<rI���o~㵎��h� n�z��-w7sӨ^�{yb��9��}��$�˘O^���F�J�#�ɂ�E�4��n�6�~�_ ���5ۿՀ:��(�,�C�M��c<>���]�
"!� ��4�½"1��C�9��-��{��+��Mn��˝�}�c�ps�L�U E�h!%ቚ��qɣ]���X�+BQ_)�C�����[�`��:00N{"�O^�dB;Wq�\���q<��Ë\�EZ���w���Wi� "�0N�R�0�&��wq!���2��� '�7঑��?k<��؄��9l#�e��a$,`�A��9���PZ]9;������ �O�R�<���,h=>{ ,<7x�  ���g��A��2y��m�T�w3~�0x9�0��l����ʸ�8��ݖ~���AO���\_]ഘ>�7���I�����P�o���!���di�ʮd�ZRI�ʖ}ɾ˾���P�.���}�$E�}b0��`��`��9��<�������+Μs��}]������>G$��v�n�,>V������Vx��'�������
��~҆��)h1�'�d�w�1�Uq?
���\Q�n&�<''���2D���=K^R�<��Ot�޿�!+���k��o)����4lF9����b��@�i��H�r��T�?���\�騊�e�8NN�TI��E���������Q�x���S�~�j̑Qg�!��k�~�u�^��~��\ �;�5t)����*u��=�%�5�?!�|��z���q���dvQ�[5�撶�Q�K�E��s%S��j��dV������]�3�߱ݳ0����u+H���-I�.��h�V�"۝��&NP����DW�'���O�D���/`)����Ǡ��n'}���<�M�<8��	����?�8J��n����vD�!��� �@jlF��F�T-^-��a�T�bF0�5��x��ӿ*��~\�o��M}��|��L$6K������;��	�e�g����w��K(9Q�z� =�E��y ��`;�����a:r���&T���En���^�����)�k�P��%�
v-(}B�'F}�G~ȟ<& �j�_j��&.�R�M�2d*G�����Ɛ�6��?}��;���>�b�_ �(3�h��^�S�8�S?>���&_���/5�W�
}�sZ�8�9��/��s)��_��_���#h�HN6�PȔ��|n2P�q���&T��`��s���NOM�U��q��٫��e�.���>X��X%�&"�^�MB�� �{6��L���%�f�\���c�ŵNOB���^B�	�����{iQ����<�l��P��_�0��T���g8�O>��T3�R��a)��}�K#�m����+��#z�����4'3	�]�-��_�t-�{����M�E,��+��e`w��un������PI��������Y��u��?�n7�U��Km����?���~�-B����<���;�~�~����R�d��q��矣R��D>�$��ŐI��FȄ�I���p��}���~y�R�tt:�t�߄5������`�	ȟ訁2�wc��+�u���$�����I����������\����c;��\ur�mi����K�+����o7�w���,���c����0��^I!��n�M�����X�O8����	~�ء��.��PH��G� _���).-qLى�5ùLo�+��Q�%c#'�#ΰ��U7�Lw��s�I�L�Lղ�����7��aǯ~��r?Q�gS�5i|?�� �}y���z_��^=��F�p�)T�6��}tz+�K�)��g/@p��i�qB���8>��	P��:���	O.��ZT����2r�5���|����+�|��_��n��4h[�u�X�ϳ�n�폙�K��t�ݒ1�꾹�[2�tM��F�� $�)�jܯI�kR��Eg|Z��B#�3�o��7q#~z�}x�w.�9�ib����>�9��I��.�b����ۖ�Kx�O�RS]��Ķ}�`d�~��yV$��IP9�r��E�{/c��p��B	��Fdo% É���P�͇��y�bɄ�=2�`U*l��3���M&y��������j����NB�.g�f���ӛ٫ObH&%ނ������j�w��ÙͽD�>O^x� #Uև�5�d��V�71u��cK�����}�Xh��x���j��{�cp'u5��k��I1��ӛTG=��;�U�!��l�l���h�{s^P�L�Z��x�Ң~��I2�� �<�L��K�k�
��j�_"�!L�����-�D��	/��Ke�>gq
�l����!�l��#��g7�:�ҾT�zs�
c�u���Hmpa�4���d��o�yo���z�i���3x���?A@�x~9u�5�3�A�&�-�H'���v��8z���u�q��_e�?,c�>���R:+"���_&!��1+�bV�4�Ժl84>�l�x�~u���.+�/M����
�u�",�R��7���\���ׇk���oN�� o��p�ƠJ(M�䦠�_ek��]�bZ�#�j�Iˣ�̧���RG����q�4�7,T��ͭ-r�~\7`Pi��%8U���;�������P��Їn�#�r��<����؃kK���N����3�,�1cz�O�s^�y��4s�%[ՍKN̯�i�rHf�R��.�����jjj*�8����Y؏O���Q?�add�j������Z�U��B�~b);S�je��٘,-��Y�b����Ӯ�f-cۃ����đ������;�]�AUN��ܼ<k��b]A;��KnW��uE�n��O��o�����L=�%�94����uxտz,����O�X���c�$ hk�W}Z��[V���8�᳷���ݞˣl�o/~���_�o:s�1B��mD�Lƹ>�-����O"�Q貲��[�T����$�;����L�Y�E���l(�5pb���E�Q��@>u���-�Q�m_iAwz����̊t��Xc��	+��%�MF^��X��f���$�4�,� � ���(yR@e?/M�����c\�w?���ɢ333&�.\���.�n�@��8�([9�W�#��#�í+N��J/����'-��M�;����SC�4��a��N n./c�끦<���ۨV$��p�ȝ6���'�~��_>����{�p'��	�&C���5�������������	Q"T�0���궕�[%/�|Ge�N��P���k���t�����-���f��ne^�N{��8���r�T�T�z�h`p�zo�X�e[�͊!Fո���g��)�pR�sXC��R��SW�j�n��K������g���L���{n�6����}�qp��*E����/�El3��ҰgO�q�5��*�w��@Q6��wv��66-�����M���k� :�G��[_i*�P6�bx)y��<���\?˻���
��)	�`���j�d=Y����Ƣ�GtI�n�4�#ܝ7J%�jp��	a����w����g����:��XJ�T�ݜ!v{�B�q~<Fqo� :�+诋��9Τe^=����h ��^�'}y�%s�A�ӊ�l�����+������s������@<�b�K��L��Z�$����D�/=(F�{�e[d��PZ潅]2ɴ���477W޶|G "��݁\!8*)9���" �4�@`3�Ck�;����sK�<PDdޛ�ٛ��B�}"Yw��T�4Ҍ��3qI���d ڨxߦ���Y�#̀�xWPP�����&�_��y�Һ��A��#�x�SL��轝�Όr=�7�i��>��Oܙ�~��hi�q���DX���`�����C��·ӈ�zr�9�+�|�x6�4��]|ZN��A��5 #��/o�]��3D���_\�4`��9�G�8�h���厝c����l�!�?''%~��=4��6�n"�dм���r�-ߕ��)|-y��W�_!X5�� G���h�z/V�ge|b��;��GA�9��V�4���oye��W���c�X#�y-�tg�$v���i�ţ���o"/7��뺁�����L-�s��k�ѣr��Hn>U/p�C6xy3����mBh t�{�o)���Қ������]��5)�V(Z1���ty7�"E�fC���p33g2�O�0ۄH���8Z��B��/�(nX*zM�~Sj�۽��H�.je����oO:ל�_r0%���u,C�1u3{1\�⏌��h{����NН���L;�G�FV* wθ��I����$��;D�Us�^-�-����/�c�7'#EeX�8��:{��9�{HH�h��I�P�bS�+!!���@�x����}ܫ|SN���FA[Ӣ[!��!ؠ��� �7-�{k�X�y����� 	?a �r�"�:݇�}��K��T����RӗJ�c��H��}cz��k����}��M�b�x���E�j�3���Vf�c �|L����ݗn[K�*gW��Oȝ[#W����R|q�Rз���q+4��}�Ri���M�6ŽU�`X!���d��D+�mM'R򔁷&��	����5���o``�D����O��+����U��Upے$��h*�5�>���p"���Y�As�N�4,�n�'��;����:ޑ~$zj���kZ�1#7#K6kA��P~ Nܿ��W�UJ�"4,��Z_��꛱�_5l��7�nN}4����$��J��q@9q+�������͛d�?�Լ8�(��"��`��|����ؼ��a
e�2S�^̧�������$n���\�B���P��X�jӕ2>ՄP�uE�Υ�o��%S&z�D�qqj"[�����;�؝NӠ�HӝDI�B�h��*U��O����D�h���*���^�܀d�Vcގ:?kmU9M�a��Wy&�|���###��u�E�nI�X�4wvi��M	Zv(��,\R�`0�!Be4T���8�������lzF���%��e���s	�	Sp�%/L��-�`E�~FӾ<��� �����0c )ZH7��M�6<nɈ�rb(�id�Y�"r�/cOʷ���O*�8��醌ע~������ﱦoRR�w��c�z���B7�R8��1o�L� �w�;a��s�؇�Ur5���ߺEl%5��"����=b��V*`FJa�-sc�b-�&�����5����&>�x=_BW��C}�<���\��HB�Fp�_�D}�=I��/��Z~�:}'bё���|�wR]	�B��� ��mZ�,%�����a�Ґ'��D*�m���OE�V�'q˸���T����\�����&��QM�����кIic�rJ���M�yyn��*'�U�\_��X%�eߊi�}��m�?����[�t@8���~o3�@QG��h.��_6��7���oRӤh�����9��8Y�aո� _�A7�ͽ^1$��p<�O�W���ƌT�����څ��&͠�W�������mT7�Kn)2�4�l�ecOx�@  ��s�vm0�����I�Ҿk��o:H��5�����6��q�@�#ťi��4`Z��n����C�%EF������G�l�l']}��d���/�U}<�����cw��������U{\M�׿�~Y_�x2,�_𔋡�K񟝝VR��ԗ4m�{Ct�7 K#��uH�n�w�`4�l�]u��M�ai�޹:M/;���r��R�����D�S�:!kW@��_ɡZ^;�|��hP,&+{��	:��/��	]����ckhc�Qѽ�݁�F�.�b6�x��
q��ЯL�v1v{W�a���#���{���G �b�PV�B��]�"��A�|Ⱥ B񺾾>��⮇m��9HA@/�xi��:�L�S���ٞ/B.gl�\��[y��	�|�i�Or��7����	$ot꺝T���jd-�=��K�K��_�� 4������K�����8�h��cb������V ��"�zc��E?� �#��v�ǞͨY�UC�������W��3�/'���7T4�yx��S%���ϧ|��<�OY�'XM��J��4�,h�Eq�,ft��f��r��=E�9��82��Tb譧��M�EfT��y�z��Еc�Oݬ=v��6�rB�6�RCzZ�]k0����^��O����g�2����6`y�]��{N}��d�����I�e���76�&9��8M\<_Y��e�ș�G��70�*7��r�Y���^����;B�@2E�L�֥�G_8�)�!�u�� ����"��ȋ�ȳ�704d�le}q�p��}5��*��:��#-�U��dH���/׶x5#�m�j��ePvp�~�^������ʞ�?_�mT���FD_�Y q�=����.pv�νRǡ�k*���qh�@��7�)'� �N �ܪc҄K�Wb<J�Rxq˵�T��\uJ��\o�=Ie{��t��U��;LL�C�KK�3���;���z{��r7~�1
V	������f�쬶��M/��C��A��Ȼ;{K�y�fu�,�(����\m��x����=��24���n�W��O��L����!���ì�����BŦ�MH�� ��aŌb��|A$X�c��AD�O�J��_�7����H6��ɣ\M����Ư���-w�g��	�J��������QqqqD�Eč3:���)" �/�KcD���ئݍBO���q��yHө�dp�����c�;�|��n�y�#'��*��<Dp�2�-2�KI����b���?�^,b� �
[ow�����Z��[g����R��Ȍ�����ʢNJ����^�j�\��[Zc`�L�_]��zY`ǘ�t�p����_g��_�z����'��r!�_�{
u�LdV��7�1&�����S�S
�������������ӯ~���y$�0A��Δt4�rl1mlQ7!��co�]ZZ�f�����Zހ�^� B
�l<ѽ̭�a�P���k?
�z��ʇރd��NN�;���mY�FCą(s��exc�����h~qQ[�ˤ[�Mn�T����g栕Uυ���o���ud�($�vk l����:�N��J@Qe��.]�|99=]W$����|���DS��Qc�hzr�D�]��hO6F��	O>�U���P&�l����8�"��⁰�0���m�,�|;���/�Z�hި,���&�ȴ���I�'@�p���>:�=�#�C? G�I7�c%aWc��)V奒v
�3ҤLI�s��}K����o�d�e��3pyW"�.�Ąy��Ӟ^^���N���8�uKM��y��������7>~��MćJ D���]���f��2�kRf!�^���� 7Mز�oda�o��P������31}Ɔc#"G��ƞ���T&9��Li�A��]l��1rk�s��j$�␬tp�2t��-�r�-e�yόx]������^F��2�PE���.��k������|ۧ����~��!{){<5N�b���^"��k��m���c��U�*�b���P���Q�-p��e�n)����K]R"��6z�7�~�k�h�`c���2���Ә���̫xh.�Ю�����%F���ݲA(1�e4���wǴĥKYfb�%%%��f� 8��(.�+�V\�~ְi5�E��-M�p���z��r7T�0����q�32�w�,,��A�>�k"�팩���'8=5E��K�SwvG�t�ŮG�.�Wpx1ܯ�lV����"UN�Cr�����;Z�)~�����Tn���f
�~:�pϦ��>�@�x�"���8��A�'��,s�������_��-^��-������ew�'�O��=J�el��/�a�(g�;��7]%����1޸Rw]��E���&2��E޵¶
	=�1X�R����������e�C��#x+G��k>3�$9m� {�����ON�T[������~�S�tjj*�O������/�>l�b���|)��^sQE��Ǹ �ݑ���vz��!�[:�bb8T��������[�I!����r<�WUIzz{��.d�(��I��c�^�1��ֳɟ
�<y��qc�Tp]���Znq���1z ���O�Aؑ%DО J"�nl�w2��DӄF��@��w-Y�!*������[90��{s\Z�͆��� C���*�;=/)�D������E�5P��=h��q q�ҋ�"���~t��!�D���M)�x /doo�V�@�.r< �Y�W���!^����5����e��_�Z�O��w������{��t�ݛ�v�-�!J��!1a�����ўW��A���� gY��J�Wm\_�}�8�����`uӕ�e��l��r��j��L��.h�Z��D��f��v��t�q�6�G�*��D���؆w�l���C��/�k�.�~hȤ��"=���O�&�iԛ6���x#>�����+T����y��D��ŷ��Y&�<А��^�l������^����U��cR��|Qi���0U��� ��wd!*�Ǿp .�����:Q�L ��M�g�oVZ.,�d
�P?%m5��K�3�y����0�qؙ�V�9r�3����0�JgQ_^^~�~�X����is��n:��N��R6�PP�g	�/��Y��MNN�]_�8K�+(B�E�h���7���x����*�2m�sxe�����!��$w��mn|�uϘ�M(�;�D,W'�� �@zY[��_�wN���@�9��z�Ys��EDp�))����Q �� �Lh.�]%��.�q�
�=SPÔj�C�����}��BPCׯzC����ʰ�:�S�P�� �M4�G	���W�a� 镍��|zS�6����%E/^���˻��LMyO7�m==tTF=�&��ާ{�ӂ���^F5|�c�����4Q�.���tQQ�d��a���π��|`��ge@���t5��O��ry�;p ^D�Z �����v��6@6��2ǡ�n�:�2H$ve���uPI0���
{�1ީ �Ey�;��񩈨����T!C�Y�+)u �j���X:O��1��0�}Y�H��V[�����n��E�ʟ�t�U6�4����
s'�o~yYW����8�xc���##==nD�)ej��Y� O����@u������[��;J���Y���s�������%�&o��ء~Wf��}c<ژV��ck;���`�(D/��잞{@��׹$5��N���-r�L~��D^��f^?�i�i�A��)\=��!�]��n��qv��w `���!�sXl����s���lK�Y�Ԉv(��
{�O� �oiъ�^z�Jx�[�#�|P3o���jD�S���bccc�蛪]�s5��!�����A�4���S�yvpyY����!�ur���|t���IA����<ѐ�m�����F�����B�J�?(%��H�ಗa>�)�*��}4bz%�F`���q��rt$�27��v/).^�tn��@n��~��n���NkG ���n��?T�5+^A6QW��x���g��y�ƀs�ZG�Z�w�� ���q#;B�s���4r���� �e6�[
x�����X��M�P!����;��ixZ��7/��)^�O�vk��z^�Y��������/ ���1�+�V~D������C��ɹ�S\����c��tG�����s��/H>`aq�X``೨��7�7��w-A�q��V������ ����%�j�4���d� ����ghNQ镴.����J��8Hu�aN�� -|��@o�]�%�!JJ�ƒ/d#6�q��/��wou�^�Tx�lS����=��R'����� ���s�	H��#LL�u�l�	�'Bx�,Z3��<��f��v����I$��A�S�	1Kߡ�%��@��k؇��E�1Л{���sb|�L��� �A�o*jk?���| �ťT�c�ةO�Ү/w�L�q(ѫ{�iy���nO %�OI�� 7Ź��c��!���&Y�L[@��*�;a�tl�N��A�ɞ#���r����)�V4'�<Z�p!B)����K�f���F{''b��\�
��-/��PP��(4P�m/i�)P�P.���Ǌ󤧹SҐ5��mT�:�b��\��~I[D��~8��,���,��F3PL�%���.EX%�coŋ���W:q��0E�T#���S
4{��/䵪׼=��9(���$A
I�UO!��J�i8xx|\,<��t�(@��b���C�"����&O���}��50$3J�,op����@���ֵ�Ѧ&�<��2ẉ�Z����t�13`t�W�Hũ�����Cddd
������\�)�|9�9����1h������^���� �9�PX�xɋ*����v��vU�p�36�ܰ`��nKHHȩ�[�	t�P��K� 7�!}6~��ThEI�n޼��cz�~pFt�V���nB�h����_���(Ͻ�<IR~��8(�|����f`�������i:D�wo���䲒sq%����\ƞ��sAc���i������\D|��{���8�K�ƞ���\;����Ob|?-����i���҇]o�x�>l=��az[�B��.���xs_?ߝ�}G�e�[��Q|��w�+���w@�ކ��)���	��0�\G9�'mK9��|����~�	p0
p1�䨼�z^=�*���ɐ��K�L�Jq'�o�\�)T:Z0�F�3������Ŗ}�X����-5��=e� HUw�`��͛)MMʴ|�(�?G�~UN���D+�I��aB�<iD�8G����2 *hOEI�400�O1��Ki�L���Z-R�S_�~G�5(T��rrr�W� ��w��%̨U�`���]�.���l��˴���g���jM��g��Ѧ�����_���R+`��K�y'n���O6��4�E�X�:��x��ld`Z�!!!��Â�G.+(ht��f9S�U�d:R��������yy�v(	u��:Ͼhn��՜k�+!�QP�,Z��O&�[�>⤣�$|}�o���m0�������b�i@�-��j|�e���T��0������$��/������g~;~o	Zq����c�}JqG_<���Հް�٘&0�V�8�bu�W��G�z������V��@|ow�߀J��uB����:)���?c&���mnn��I�(#�J��ٿ���ټ�ѧ��ӓ���pd��U��S:�3f3��C��n���L��MBB❶�|_\)�Х�h�(���6�����(yo�q�	N���h�.R�&B�t�͟��?6�;{�l2 <ކ�v�@����S��WF#����JE�m�V3	�4�x69�=1a��fϕ�kL풀񯮮�V[>L����Py�2�\��:���L��{��j���V��W��o1�T����~�t��yb=����,JS:�	���M��K
�G>���?Z�`5P�s��t���i��۩���?�x��B��%T�W[���g3-h��3ʚ(e�?���ld����#��ņW�^�sE7��D��'���G�����vZ^��I�1d�8	%�Rb�B�e����2~o9���`c�&�z�R�ġ��bZG� h�{�H���g�&#�ֱ2��i|@�pf�j˶���a��]�i>r%ee�Ui��&���-��^Z��2�-�~aZ�l�c*%ݵ6Y�XU5�.XڀKv(�� �,��@h���3E
i�t�����������?���@ ��(r�g�_k@���;9�,��ө�<f�=��03�i���􅬍|��5ȣx�y�6J����G[?m�|7�l��$p�LV�Ł�)�aXxNǱ�R�4�.3Te�Sq}Z���~���Zx�,�-8�^�~�P�gRISmIG#�+/S0B��hD�̶����9� �Z��m����G�ITە־[]j��Q���{�׮��v���ԕ�ѻ�$'4b�7
W�Ҽ��$gLU܏w��\�a'�ߏ"HHJ��8#^�[b4�V��-6���Q޻�ߌ����*ǡ�H�y�;U�e��o���q4�n������ݘt�"	�yT���C�S��\��}���l�}��{t���ͅm��i=Gtw8�y��=ȴ+�Rc>��J�����x���#�wrv9�s����gU14y �ѥ���Bj��oı���Jǵ���<��� ���9w�<i��D�
'Caaa��������v��r��.���T`�ƕ73�y��i	u���o������C#,Nk�k]xg&�_�p��y:����bQR�e,�R�#R#�91��4!?w�r�|Cãq5���9uuuh�W}�^����?�����Յ/H@��F���E���uA_Hw�bc�nς�f���gH���0��/�[%ԁ�D��TM׉�HA�=%�n��`���`>*)3����e�HN�����������
x*��2w(��Rc-?Z�h ���S�黾zU�0��11F(�7!�o��)�Nd��fޅ��
���w@��,/ȣ���&ct@�m>	9���"q��h�2��_�:�	v��+Wtz�.vv���f����<�H���RM��898���J\�}[��⌡�˷�a�u� ���V� �ҩS-bo}�� �u�.s�֌�+6e|N�`��ÄW��fbZ�Fa߽r&�������b�7t��������aȵL�Y�L>����ձg�}����v�4	p'���EP���"�&S2�zG3#h{��W[J��lii����r�����}K�jM��  ��@�p�w��)�W���7lQ��v(@�4�U&��� YlG�0�����G�/7����
>o�v�Ci|e��zp���� M�r�<�z����P�����u�@���HM��v�=zSp�F�=|Í������ �@�p�T�U�_v�#A�om��ҏh_lT{?���z.g??�p�׍tٕ�:P�9 ��T��nad�U>q�C��Y�i�C������^_��m��Hˣ~a��1�=�Ҧ�B&.�Smn����oRS���3ihi#��L�*�ܡ{��������u�7�N* ���^��D/�����������֣����`(P�1�}��[�&������?z`��|��*�0���пvܤ���z��:���.%���.<gn��&�Mw.���c���z�5S�}/Χ�Ӕ�PFg�br�-Z666K�KKW��8����ϟ��o� բ�c�;`Jt�8�m/��M�>����cT0:%=}PM�񝞉��h�ʓ B
��[:48�4�!�$3��\ -j�4\yu�ݫ~0^�&��նP� ��Ÿ���~6SŧY=,w2,Y��<�6 LT%;�Z�B�R���Xy�1�=��dO����S�e���S�B=_��t@� ��Sox�X+�1@���VQ>nNQ��7��JUϧ�g�o�M�,_L��
_<��i��'�
ڈ�8>>~U�|��X\���f�����&�t�y�/6��}�c��\^� r�����{i����� ZЌ䥤��I����^KŦ�&�R=���{Z�_&���&d��� ���)�<�Ī���:w �d�Ps�s@��B�j[��I��!�	ך�*�'�����Qr+q���E�������X�Ƨ
PҠ�9M��_`7m�����y�7��MZ����K-�4#^GRu���LY�ٛ�f9ݐ�*+���xwٻ��(xK���+�:��\g���%��WvP�3�x����E�G�l����[��3� �1�k6�nᒎ�2u�tW]�2CV��+�������K��>p8��2o�C�C�95��Q�r�i\[���,���0���i��� ��C��\�1�l�9���K��ɨq��#-ҋC�cz���}AW&�����կ��&_��S�d���Ҽ�&�o���ή����6���Vɹe���[�U�{|��5��ds��v��L�e�s& S�zՀ 5����p�Cbz���&&������!JJ �O����~�q&���b����G��`�xs��!�� ��t7Wz��B��`�m<���~�$4f?�-���ɸz�N�+��K���j%��s��_��ݾTt�z���' ��EZ�,,�&l�A} ���_ s	O�1t����KR::;��O544�������Y ������ɩ��[4M���J����?@L����`l��#LH�����Ƽ|i��Yq�Óϙ���Y��$�0�+����v"���ƆL�$+�\9�S���؝)J����� O�V���J5�Q��׼�O?�C���SDw����-���*,.V���8Ӫ�_;��k{9�����vQ��N^8��� R
�O�UW�+k�鳌���?rRҖ0�9���`"�FGU;J�M�t�GLR�#Wkԕ��l��������X�y/�.����%A���[
/�,��-���+2v�j*l=҉P���14��ɩ5���{X>(ܿ���KkF9� ����wr��
�r���ݏN�(9��tߙ�`��� �{/lXe;כæ��������>mCCL�)pQ#�!��
Ͷ���:�B�o}��W��r�c�F}���ק�]��_��wtp��4Y����t��ͪ��Z�U��UVV^�b?�D�Nk+?iF���&�x'�ȑNk��㘪+���  �@��:��O[�i?(%_����ǲ]_�r:�J�ȼ9M؊��=8*�!@3�s?����nY��|g�&�JLVU�Fj�(��L�n>�B��d�X�����c��ԑ-5���� ^���[[�,оx�$��&���i䱦�b��. �wYm*������ ^�z@>�M��1)l�f�쾂p�
z�����?�۸�B�E�4$7`&���j|G�k��L)����A�gg����;�w{�$����rr�&7//�6���س�4�o'�mf@&<8��H��CgI��0/B;�.�>�'w��q�>�cXc�|~���?�T	��n������'K��(W�ِ��g�On^͈�rn���C{�`~�=ei.�rZ�C3�@O��`Y�h�#���Bx~ء��K
��웞g���)��4h��T��*�@Z(d5�������������Nȕ"�^������ni��>����j� �\�o�(��i"��7>�z����-?ڵPOY�Ӥ���� R-)9��,��cm���]�����i�hj膢"����#%�fɂ@�m[w���уX-�]��K�n�v�iT�OaKspd��+?���l(D9���ч���{�
򝾐d�Ԡ�X��;%N���q=]�2���w>5zv�������O�
���1�'~c��靉��;5΄(��h��'�����{�)u��� IZ�t�ֳ/�*1z1����_���s�%�A�GW9a��]���"�����X��о��"%4���c����Ug
�d�F�X8��ٳl�l�? _�	\�'���¶T&����M2jj2��^�Ue��S��]m����y��wX,�*V8�`q��6\����\@��+�q�s����Yޢ��?]LH;����醫�]z80�w�E�Y����1/�?&���?���¼�ؼc�"~�oO�{��Ͱ'�SSS���z��
~�ѷ"�ۃ���ll�L�ʧX�'[#;�i���́m���2�tG�/�WSy"Z����I'LՒ��]��I2e��[KE�rV�p�0SQu��d���sl��1QQv�C�Ug����z�= À�&C��ؿ�HVm<8B�@��6p��ޅ<{���y a�� �����Su\Q�Y��C��\�J��s�&u[A<
^�m��2���5������V+_D���8p�OeQ11X�.�ح�l����L������)==�Ψ���{�@$X�l�5b_: 4�ᶓ *|�N���p'!�.��Mz�OB����k�x���DQ|��\�fI�R RZ~��Y��Z���Z�l�ߘ��-�!�D[ ��L<��Km����S3��w���Rƾ*�!.�����?���F��m#��d��H���"}��,� � ���c;����v�oSn����������X��'�(��A����]�o"��?��y��ΜZ����m{g�_���^���C� (ȸ�rF�OF�b�u�����w�����ӏ=6փ��l�8��!u�7���o��4�&Vt]]H{�6%���焉�e�����g�΅����3���^�H�W�H�uj��|�<dj�!R������s�L[c �Z�,�b�X�#�ZUŵ}��R.p1���'�m��u�3��w�uI���iۏ,�g�P7e���[��z;q�ٺ�C��(�1�pzH1*å�w3MHx�s��	D�`YWA�y���ӎ�d�$�����zw�bTt����P��4t=�dp��%�l�.�DaΨ��jﮩ~0���f
�!�BBR���H�[��o-�(�o%Aqy���m��+��O�w�H�������fL��zL���20>�o��|��/Y`��|�P��0�����Z��f��{?aj!��۷��AL:n�	��4a\͌ �l�����Ù�9_�_&�O4Tч��(��q!�P�������\0>{(�������d���9)(�88/���#��'�9�%BB;E�Hh�Ǵ�:�q_0��{���nw=Oq �4���a�	�(������wҟ?.�!~v�w�|���9�]��Ib|~��:T������U�(5���3r뒞b�v�HBE�ty�^h��e��v>%^p_~��}��T�TU���C��ͥ���TWY>UMy��&�.~� B��)-��w��_B��[}��w�J� SqE��YZC=�B�J�R���*�^�� �@�y~i�f``  ��'N�|��ܽ6Ut)��ʧ�=1A����:D�k��v�>�7�hO+LD��E�|6�cpg8;=?����x�>���?t9lK�O"��6��}z#{𶔂B	�l#����Kޞ�v��� K��Ъ �ot���r´��ў���-���/�3g�m�zz�FG3?��I����������.Kоw��-\������%4��yk��\9#�uf��MP���[+eu6;����d"����Yh?����
��Ҕ7o�o�Y�'�2�&P����b�ofr�����g�ܴ��M�K'�.%Yd��B������}&�98X��m(D��B�۽�w��ʉ#�K��h�9�cP��E��%��'���w�/����y��'0���\�%ȝ;z`��ʇOq�b9&�e8����&���Ie������u�T�ZX�]���~>P��߇�� �����4�Ml��t�srptǝS-t���
hzs;��UFSUԛq��#��obl��t��7\��A7�%��1�a���='_�sv7�53r��Fi�P8�B �c�9�uu!���Sw�Hus���m�m�3�X�$c�
~���[u$dg�����q��˹ߊ�z_����S�ůƕ��b�k����A��V���,:`Z� ��GO�C'��>��V����
��M �;TU]�����Ӎ9΋,��7�I�n9~|� ڠ�騫�qm�-�'�*�����e�?��*��uC�JC�@�Ll7��(�9
`����ō��~=��(4�F>����:��Z3��HeM�cX�D˥�=��ڎ�@����?���8ύ�y(�.�R�5
&7>��j����z@e)&9p����� `\aE�b�i˄L`�6�ٳ��
�����:Ҙ?\���v ���Et$8��Kg݌�~<��"����6kQ���c�Å�bWVW���Us��)++�t�F�R3�r�������Ri�d@�@�[���E���q�w�#�4�p�r�D����!G]p �ju������c�ys~�fV����/@q��eb�ImR��.�Z�I�Xx�����D�Ϲ�c�{	P1�W2Bg'�m����l`p0���CI� KBX��KDb����n\0�
����!���&>]�5w�ǘ�
�g^tc��7��K�˲�EJ��b*�S���3���iw^�y�ҸO��g�Bش�!��d�3�Zr<�%׿��#����#u�߾s�@,����O������#�`�-Y(��ɱ�� t�~�n�ف������ 3��rޣ����i:��ՏGʁ	6�R/Q�	AVz�E�qoO��G���bޝqZ�90Wy{x��LEmFo�1q���;`LI�C��0Ţ�E��J�P:n�Sȁ�zo��O�7�b�:z�9@4n��+��E�8�Ή���쒐�)�����W;��l�B{��$��=:�L��J��Ó��l*  n'"���<S\��d���.l�n�#QOh6�c:�@UR�	G��>��3@�	���94�2�A�yǽq�o�_���2c<}M}I��d���T���5�Ǖ$�	|��r��cWii+��:�t��+��b�l��R��'����s��\�t�j'����os��M쌕�"+��^G�gώ3e����=#�\��z�(�/~tEDR	i:�[�i�$��Ar$%��C@��F��a�����|��<�y��c0��'�^{���.�+�n6,��H�&<`���ef���%�g8���e���·���U��VVy��9��٫Y�ж�$$nBi߿k ]:��i>ٟz��I������ǒ����&���"���t�_���������B�;��6��iأy�q�(��/V��N��L���`���6��2�wq%�f[���b8PVM�ke�>��qf�(#ro֛���8-�av �=���{M����Z>������AL��r����b��$b����!�΢���[��P�^6�I��0H��Q����j�eG±�:�>3?�,��3�;����h����[���D��/]�Z��Um���O�j�':�f8����߮�lo��͗x�*A�F>�Cm�BW\��p{������ P�������k�NcK1R����@�kHX��~A�9����=��� ������2�n����C�͘gG��_�˫����(�P'^�h���T��m�C�
0�8���%�Z�B[A�!"�=�D���B�x"@P�q̖����J:ٺx츂��B����X#tycV^&F�䠬֍�!�S�;��GYYY��� �ҷ�2����*'-���2I����>:4c+`�L�	AvN���i7��_�k֧�9u?�_������l��Y��W�vy��8��QOOOB�e����0�ttt��ɗ<8�o�LLȞ��
X�1Ǫ���8<~��ߥ���'t�b�z����z��� �}P����u�24��2�!� `�v�̽�<wRQ9v�7\Qp7��?Q	���R�Ӝ��'�!))�5U|��Ho��4��@cr��:�-c|
t�ҐG$]ݟ�H.�?)ᷮp�;!S���=*nmƅ�}]i�x����Ŕ��w+����%��n:P��G�ˍM��c߾E��F��Ӫ�d���r�ZҺ�Z�Z����	�U�����C�ŁT�@�%XH�/ޮ��;�M�r���y���
aT�:}�W�а�"��ma�I�2?\]�,,, !BA�P���Ȁ�	P�@�IH&�A��n"ns���F�A�I�x�ӵ1(p�9��i���W�uq�OWm��9V��!��Rjv���r��)@U�x�,@(���\�mp�8�����@����oܳ�?<�fq�@ �K�2v��'�N+��^�\Q��*oK&�Vne��ayeY\�����go���|^ʈ��y��N�-�d��Y�\诲�[��.���M��?����и�q$�v��#?I�db��c(;zF/%�gWQA�z
���L���{g�ūW����ݞ�k[[�Rd���9��ʫ�)V��~Z����;:3�������Ά�����O4�����n�"�+�m����u2���W�*�m�O�	������L4���;�[��|f�-4��p�2�صc�j�ʪ��wPG�,�ƀ�4	�C���} o�Y���^r�����L_Fu�{����.=O_?c�U���n���K{Ճv��Z��X�4�_R���U���d%�wQ��_?���s�D�QZ�3.�"��No��OΜ�<��|21S�L��Z�_/�ܝP6��XH�`ך*F�����i^�
B�A�,=�����7>&�vZ�V��*�^��h�PL�-�bmN�M���?���DEE���{�c���T���[�e]�IQ�J�zx@�1gxX�1��[�,�OAR��uA�+�,�h0�L��h�S�Q��<�Qr*�W�F�w8��<#�R?�8]�zR!�����[�)�� ��[s���v���8��qQ���O��N��#�i�ݻ��Je�����߽3�@�JP8W�!�[��M8N/:<<LP) ������L���&x���^=��^���M�̿��$"2Yu��Ą�Y��?��}z�Ҁ�l���������zӝ1��UW�H�z0���$���l���/�=Ugo��Q����ý��|֗'҂�יVq�Eݟ�3�-6���PG����1�~��Ղ$����w���mRv2���]!��)ᇐ�P��*
�!"R�ק|�uNbb������b 	��V��t�v��=�qLW����Cer�jQ��			QO�
8))�T�i�5��ڕԶ[`U��9)e���mL�@/,|8��C�n;B�B�QN��2],��Y莁�09�)AMGW`���f'��i�,{{�	�F���ޜ�Z$Hm���z;�b������J�=!�p����DHd�'�j���Ƶ�H��.�{��Z@�c�'r�ʁk�Z��: V��҂כn]t��;v�p����}��iɣ�N=r�O��_/@����S��'W1-���E	��C�e�9�dw���cE�ڀ#ϓ��ӲʃW��������d=���J���|�攼&�^�M߬A��Ȉ־�
1�B�UTp= �2Q�Se���ٍ�:�G&��+C��:*�?l`��V�Nqsuz�Ҳ�����D�o��ma\E���*��8Pr�e�	���ee�E��MMM_����A��<��QE������zӋ� �!~ʗ�[��!��RP-@�
�]�"�ݩ��V��).�����}���
$Su��;+5���y�pO�S�W/�tcj���Q%����nEe�ʏ���r'���ԣ���>��S�^o�^!��o<?s�y��f�>��?�O�PQF�L��������I�Pхnո.��}���B����F	�>Y��	��' o|߷��}{�!��٢���3n��������.;Ŝ�OԜ>/��h��Ԕ��߳�O3����y�ECb'�,��6��K����a`����ʶ5�4�nX2�su���O�\�����즋�/��9���־�l��_��݀��f���v���3#{t�ՍK��	�t�̇ք�_3�RT�'@:�F8�e�Yߖ)l�XR����V�vHVx�zS���O{�0�o� ��L�U��,hSB!z���qe��I*���:}�Y�����D����3�!�\�w��^:w���y��!�oʕ����><�Ndqe���T����Y�ʐx'�<lg�Y8�y{YӺ�~�rm��LW�Z���[�c;}D�K]2w@���"�ݫ��qA�y~�	�"ɖ5X?����B���7#�˫[�c��}�:�ThKw"yV|��&lޝ����痛P˗Zy�j�\��X��/�S?Zr[�m����8Pkk���B��T�^���ꂧ�v�~��EI&�o܍�N��K��6�
M�<T/l�������b������r��I�z2}���߽�����J-�X���ez��@��j�" �
eîk��uEÇQ�II��֯G��ĉ5�8&
�ٜ�D�o_=��s��2rSް��bu[���@�O�e(h&ȜӒ�5���Vh_D���<�=�΁U##G�ʊ�%I�����	=�b�o�7|��[��J��¹;�}��Fq�5X;���O�Uu�}>g���|��ŭS`T�`ޑ��y45�cJ�-`�C	ؓ�$��:�"���^@M�z�� )?�Ѣ7���P�-5%�����~�_�� U�y���_z��ﵜ.�PeHeJ�����A�iO^x�e��'�����]8ɶI%�,+������p,�:a�H�>nJ�zF*CC[�����k��c^h����j�'�l�f[s���u,���:�&�P�5C6w�O&�z}[x�[��?78�\����}"sOU�:�)_�8k��#�`�>�u��3ޢ��V�̃;��y{��{Uhܸ�a�a�9�I��q"\���<WP��0��w����U�U)E�S��Ӂ�����ޥ�-:X6��8��CH�c{�N?�,��:��YTG
tb}F�7d���I�Dc�9l�0�F���yx���."�;6ړ矿�j,1H���������m�H�H
m@H�i@�B��ʚp��.iC�(�,I���M/���qGVx�KdZ����W�����9@���]���+f)���U�,���DB�\�!o�Q��{�wa����t�E�"�-�<$i��1�+Tq:��]hKJURc綜V��ֈԚ�&7�G������Kx��mI'�~/	N�F+Ey��䒙���2��m��j|�����W1��
Ub�bQ4���s-Yw/��k�, Iae�r
tG�Ǝ:�I�@�h�ԛ�~�x�Y�j} 8���2��WTĕ����w�6�H��W�
�����i���['�yA�,��D��ϖFK��j~�&���Qﾫ�_�7666��׳:Yk�Gf�H��/��w�s��I���	�z/%�50�+�b����{MNy��"A��6  C���QH�i+z��a�.�b=A�Y]�Y^su@h.���BW���P=�c�Q	�N\:�Z!Fb��:v�
�1E9a~�\5�y%8����9�G7h�g�?�jb�^P�d�����Hu��5��Eِ���_�v���$�.��"Zh���gUKt��xF�j���-<+/-u?�m��^��{h�j�Ĕ��kӚ�&Z&[SB�wvv��{�����i#�5����]hߘ�>�G)��܉pz�iQ���*��%������'�
x��Ej���B�g}0tM{�ص���Z��D�]}���">h4�^YY�qq�y��L��ǣ>�89�v//����P������j�o�22
���� � HH\JB����d�����i5S4��(!���sr�*5X���7.#���/j�q�YNA�]���U�v��E�[5EyK�����)�1U74��bd��D|ŵ1���]���iճr�UPئY�[\0Xj(����%��b4m�mS���_�mm�V����YD�e��&�U�H^�- q�����yq9���J���?`�]N2e��=��u�hҼ�JA���]P����M��;>4��:� �<�M�.~rr�����4j�Zu&�ۤQ���{��h�NG�t0t �:��ODc�dC��6Q@���]/�z�����-�8�������nW���g���YKC8˘�އ��dw��� ��sN���I�g%Z5D:K䑉QF�$�e/�Ñ���W.����OA��VTac���K���g,?��9�n�^�W&�(X��KYt?��Am/�}Q11B'<�1��]p���~�T�m�t��k���$H2�^��D0�r��}��~}{��&laڤ��f�*���������Pn�xb����V�^��\[ul��qQw�����Z���뾻�"n=����Ľ?`���I���j�]er��^�Cs�eR�T�0��h����]Y�6� , ���'Y��yB�.�@���
�u��o�3���؇4�,��L���wQ=;��S2�;*�!ɭ�D�NQ�?9���(�ڪST�(��g�#õ�v�:5z{�>�t5#W�[��f}X
P�@��Bqk[[Nks ֫���q����`��1����,Ho߿�0�Dv��[�@1��b��Iܨ4�6��t���&/�\���z���K^���٩�<
��8oV�x���R��]��u�W�b[3�]aQ6��1���M{�XI	�}Ļ6�� ;����\�.&�Gj���<���@Dt\eeL�Ie��p���8-����V��A�H�,�Ȱ������=��>v�(9TRR��יn����A>�y�u����W�V
� ������6o�ԅ4Xr�٬$tb���y��Z0��t��i�����������زM��,���.�/��6�D���������|��Ne�2����B����*p%�ׄ����8O*svͦ�/HKl)�5w V���Bނ���uuM[��޽�P��+(�+�&��C[�����֞�t�Φ�����
,�E�ք�L�R>j�Z?�?>����:�������K�Z�P��J1جƅ́���m���M��3H�q����I�?���8WP�h�����C*�clzxɘ*��1��u���� ��XVV�7o���5��)�1��/��?K�x4ϖ���<��V����9� �~�Z���mv���|g4}���~"���u?_ߗ�^��K2< �J�T���d⿂6�그�^�
�!�i��

Ớ���ͭB� m!h��~}�.�u"��yt��%�B�Nx\����&@M�O.]�cf�l��	!(h�� !%�k�C�$�XAɺ�y�9'Y�TM�_.�5�7iHf���f=-a�Z_޽?׌�\���W�kH!.TF�F�1�F�j�(:p�m��xuZ���q������
�����2��%���I�WP� \�v|�C�M����3.���		9���|%V��)�*B@@^h��M�m~^�G�<�Y������[,��C0�+@n"��MY�$�Ϭ��G�9�����s�L�F=_uޥu/.yP��-�����z>:��!$z]�ׅj�^ > K�%�>�F��
��S�|��kɃ��M���ad��K/1�:�âDu�n�on�0F{���F��&%K�^i��a�J�Ir� ,����l�S���(Z�|z�IiO���$�F[��p-*Y^~P��m7{~^���f)��X�����oNr���Ub�N�YJ�V���l(�����]8$3Į�� � bݽ��f���񡦥�7�RLQ멱h��{�
�.�qP���l[�ˀ���_�Hޏ����{,0�X6(G=�Ŵ���l�ymLTcv�6��,��˙���y�`�º��u ��Y��S��iZN..�Z:Z`�D3
+**^�[^y)�?a�Z9�	��������`%��$�6}	�)��h�M92-����^��ʴ��4�d_%f�>�Ara�е�#w~�F�	��B�
��v1;l��rH���1�s�^0��D��+�-��F��8�J��h�ài�~�����.��#��ad�~�Q6��O��:��4�Ǥ�k�]� ��>�;S�֓#Vih��9t t��A3�vl�ׅܥ$xx~���9��(ǝ��O�M��I����IfUn�R�� �Ϊ���(r�#��H��v����d{PP�2���M�}��0�~�@c���,9���R�;��	�}"�!��2mS�|���_�'�&�sn��^g0�Q�i���h���e�}*tA��N�u�`ܟ�^Z��7c�S��va/W��T	Ph ��,��v�0ښ	��F)��eb�J�~|_/�e5�.v�{Jd�u:Ql<�"��i�RZ:t��Aɣ�%��\�02�B%�BJllp|:��@=���67�V(���k=\+�&��r�a���$�k���#�G7N� �#%%rZ@�٫1/I>>W��G�ߛ)�\���6X,�ڙ��g��,Y�EMC�����%���.���c�KK�o�}�z�y	���	���a!���T�B^����M��D�m�eNj*�0N��c*q�k�	Mxy�U&�^]����@�T�se��K(�1���1�x���T�7h=1Ԕ��=�Y*��+&[;������v��%" ��h��l I�F=�C`t���D!�]�!�����}������K/��L��b��� � �eJ����ވ�@u��w���-~����l)��&a`�6��i$�ͻ����,ߗ��r��RA�I.Ԙb��eZ���Gm�4�L���
z�0�� -�j� �
wQ�ʶÇ�W���#�[�݉���Z���4��7�qֶ�����8�\�b]m���i����@%eݝ��(�UF��A5fm����Oݍ�ٽu���-�l.�hj+-���\a���ѫ��}(^Zj�'������A�b��?	u�)�s�d����6Pe��g����Iq�"¯_�m��<=� ����:����x���CΈ��V�����(�m�P���&F���*4U ��Ҿ��TUUE��v�hd��CݍXU���
�f�I�8�����M���4ť*���Y�܄\��B:Y@���G�� ?s���L�?�X��RHhi�@ĕ���TyF\�/��Z�I� �Qf���7���47��t77#��~΁�>�~b���D�������Ww��"��!��ʉ���Nʾ~%�*n�{>�0;��C� ����YZaA.����8��E~=/�����GFF�Jzaf,�h[�נ݆W�MG@'�+�R6޺i��Ky�6v%ͩG"5���_��!��z�l�ڽ'���a��q34s��o�������qT�P���TFM�����M7V����W��׼,-uǎ<h�ݳ�=�(P�Z����eB���$\�7`m)K��tO-��`�Od��X��$
�] :�W�-n��c�c��ݫ�,RS0��F(B�qtl�GN�.Du��LB^S)q��`.+%3)���c�hT��P������ge�|��J��L RԚ�EKlS��3tSSSs����U�5.AA�C9���0;>��bԥ.�E��!�S3T�%2z�D��;=��<Ř������܏v��3��H}\x3"֤��m�n�n����7�J�_]�����0��d��c�s2������,�F�PK�8���2)����?���Y�3�萳t�L�f�"Ham1�P��7,�ۥ6ܺQ7���9mR�����bS�a�����-�ȟ�#���Hº���N�WOrKQ��w�: �j�ųȯ�{��<��Mש����״&.�5z�l��K�׏���Q�H��G)��)��f�d&_����\]�[�t�X+���R��Ȓ��2�_Q���PC�ǚ�F����{;nz��G�J�Ê���u�_�4AU*1iyq�a�@��Ta�`����`r�sx���A��R[���T��tvz��x�%Њ��v���9��!"�F���8���>��&���}���h÷n��iO��P<����A�����@"��!ƴ��>;QȒ;�%�/���;g{�ݸH�!Rw�>J�N�<�FPsN���*|�H������(�L�M���	υS��.� 9�,ҽ%5��ͥ�i���)(0�YE���ݻ����]�Nk�*�L������FW����Pd��b�-V	��bsxD�0�~N#�)e��i/�jI���P��^I!#;����8wsn�fgg3}��_A9��N-��S�l��u������	P� į���������4�  �PK�&��jU]M-y��.���ܨ�T��]��3w��ͱ�&eCcJ^��������^A�Iu�al���!���� S�N��s �Rr�'9���hպ�u�v�r�n���Oܴ��[��¸ğ�@	�<��q&�҃��e)�k����(t���y_�]W�t^���{�n�r��U-.斜��6ض�z�d<N����e+�."]]�U��Ҁ��ZyEP���Fxz1ꨋ�9C��5'/A:�`�gr$��^m;�k���Rlw����*d�ЦA3�u^?�ym�o6L+��:�*���;�6�clq�֯_<�I$~d
�C5k�.1���$ �5\"��X���Jz�	�JJz���'A����:G/	;Uy�<h��Xp*����x���z]�sYu���]r����	�,Dq�^6�9���0���u�4�w��*X_>O9�&|L$/� ���Qh]r��bm���\E���|0v)_[[{t�/~�v������w��������K�*�DgM��M[�Dt������Xþ��Љ��3�7FM�SS����ᦏ���\}ɫ�D�sۛ����4ৈ�s^��6jp&����o�5�4���)u��X]2H���(��0�����i�����w|)j�.�@ˣ�z^V�Z@�[�s٩"o��<�_/ ���3���wJ�}��{���p����[NT	�c�
�g� �>�֟�����޷�dR�!9��غ�9\.��1��)|,I)���c ߁���h�I�`�|��<����n�,"Wi���}�q�Ag�X�0&��O����RG)���졹������ɶj�5�����әp+�_V�@B�m�&I��'a.T�ot���'�������(^ �k>|x�5��ȯ_��΀��Z�6�����*��T�%;?*wu;?6�5X����+�公*�.�w/�NMM������PGQ:���K)�n�w�o��D��@�<Z]��8GÅn�4����{���u^�@<�$k��xDLY��H�ˤ�W��76.HII)��D��)t�Lm+(00ӱq��z�Cc��#����▨{�)v��>�IQ�XG�O� �W w���za=]����l���� `B�,XNN�ፍ3�+�^[�mm����� 5���4��q]���V��;L�|(l)�Z�$C��=tyR�c虂��Uxn?~♜ @@ñ��]�&x�R��>Z�\�����Gu��WK��k��s�G��OM=���ݱH賴��}Ʋ$��y�w�T�1�K}_1:9p��2ь�R�G|��ܾ>��z��f9�G���,�׮]��#{2�!���+,\٬$�����bbzO�����f��ʄ���o�j��Z]��)]�c��y��*���[��5u�⫚���&2iJJJj���� jH)���)�Cx��t�A}J|�S�ĨB�5�*�&�.�,ӞR�i��M)-�<;�6Ԁ�p��� w�N�#�yR�a��v(�P�L��`/Lgڼ�����т�6�b=tNY��߫/��^�kx��;i���^C���.�����O�'|)��54����� Gq���X�0��T�� ^(,�F�w�:���[60>�����Z�#��L�Lt|~~>~�b��:t恺٩+q����oz:��	֝N�9{�U;�)@~cO�k"��5P(�@�tSp9W�	�E$tU̢��������R;Urguh���w��=.�� �~H�N���RF��*�L���V����=#����\1/�m`��	��{X��Z�'�M�3gM�bm7�*�+�x�F_w����{����J�����#�=M�Xr�s�R]�b���烙MY���Dt�p��E����c3N�
� h��I���-�^���&�ĩ��V�INd��-�Ւ�L���p�;!!����B<ِc\%+]�X�!T�F�d�����/]ʶ�G�N�>�Ú�*c&��#(Gs������ǧ�v--31l��L<ij��A&�Œpk��uВ����aR��5A5�2��ؐ��2l�!� �VX/�@VVV ����H,Ɉ7�w��_�y�e�4h'mnp:���KHT!��3��ط0ڢ E�sv���[gS�~�@���n��~t��*�=zM�����	"Ү�A�!�����E�ZZ���("
j�?��
|n�|u���&���U�c��+ Km�`�_5�����L�~(���+J�vo9��oY�O�4W�.IP��T�0�ң�d[|����P�V���`Ogܤ�aoб�J���4�. L�	��E���}UFB}�7�C,_R�yg�w�����anWyE���sss���RA���K� %���Kt44GF�'O6^��*:H
������7��\ �<�$�3�#�ohtTg ������T���`����d�;�7<�_p�k�*��Y���<��
'�u d�	�<�8�U���C�o��;8��nw`V��͌P`�B�{��7�P|P�ӵ�(W����m�>kR���<����]�&:�p�( ��Q2´�o޼%B�zy��!��H���湭"��ḏu��;��F�PSv~�66��z�Ӌ������(L���{��G'�Jq:u|½�Wo��mV�\)��O�����upp��z蜴UԵ�kdd���ll@(P\�k�R� a���p�}�JP�~��|P�k�fTL��mU�LV Y�,�&GӞ���c	<5C�i�g7��@'�|]Ԋ���J�"��h{e��h{��_��c-�3@pLR����~�_��5�"��B"�`}k�>�/m�r�W/BA�����u�X���2wƛ�2�7�B='�c��4�>��������f��������bu��D�䉛�k�"����RR�w������}ܔ��
nm������w���4�y�뷿�OH���}�
��(�0-�!^�Ͼ��,rt�qe  L���:��T�ϓt���Y�����W�s�	����O�-nu��YW��㗉�'�Uno�k��BS+�ٱ�������n�H�C�Mhr�s�)aD�$����	:{�y�T����ח����r��H����jWWW�C��^$/TI�]dR�V�0^���ݔA��.�C.�^��#�����(�����OO���R�Z7�Xv� 햟��j�FFP�Hʬ�tQx���������B�ί��<��0�#'��N�����R���A�<a��ˈ_� ����̌z�R��ޟ�����m����_��ʭ\ֺ�IK���[[rY��;�����w+�]h	��0�sm/�_$t�:IOCÞ�Ӗ��֐݃F�4`�D���9�xm'8'��t:�����u�R���,�ǉ0(?��ŏѵ&�#5���ם�����yM?ҫ4��?i��S��UUU�DDD$������qݾ|����S\X�S��E���	4hƜww轹	��N����˘4�s�=[y9晿.Z�UR���YI~C'��D���IY�����z�<�W{]�Q}���.3�'��#P��R��X���>��[pY���kh���&W[Z�q��?�Pow�}��f��H���u�89��ۘ'��c��Qr��С��sH�)��X@o;<S堼:>ɒ��x���N�#�O�X#%.�vrr�4}�[J�Iy&]SS#��Ύ4��p���]c;<rT������-&�ئ@��H��:�s੮9^c��)ո�,��к+A�MrvVN	��杒A���ec�r\��A��0Iӫ16�4�`���K|8]��o��X�5�V��RG)�=��	����4:1�oqu��G�� c"55��C��O�%�~�Ee�<4����J�����g�w�	JLk&~d���Dia��@�F:L�I<��6D{|�r+�N��+[̕�:��@A�y(��xz�ǵ��ǯ`0l�J:���ccV�sdR�<��|��#��of��_xh��&�1�Q>�k5!	�U\��〓P��N�v����-=����3�E�Q5�?k$X_�Ծ{�f�&�-P#�����ӎ;rT�z�� S��f��:Q���}��?�����y o'z����]bbbi�,
%�"qWB@@��t������q��ڵ?���]�����t�z�f^���o�7u~�#�![-pX�����>��0[Vb�鈨����|�6I^�g}ZF����^3�X�'%���%?���@;�Z&��%%�<�y"V��!���F -�-���'�#Y&���q�t5�=_֠��̌��k�tb�ٌF�r��K�p���8��Fbq�kpڲkc�KO2��n�����;��1WR^�b�s����s~~~�,4Q��6�k�@%�IB9�Gջ����e��:�΃ާ�&HO.���
ї��,�O�Qq}�Q�磞��n���k�o�v-�Wb�4���鎂���5c��Ҭf���Sw3 ڮ�9 �	�r8���+J�t����������?���51����<.��T�hc�25��w����rp*kR(� _��	�L�;R3�k�ɫ�u��g��22U߳���*)�L �����a+F��~Cߦ�\c�D�~�5CC�?j�!5'�>��@背�{�Ne������_�:�;����jIQQQJ۞!�^�1�`P����?yʡ�!��C���ˤ�66f(�������'���75�A���Rj���k��>ibk
���%�3SO�:���X�dni�	���K�=@�n4ʃ8���M��}ZM��t�}[)�Qک���:��"�V�S (��q&x�h����<�Ǳa�u�\������m��lQ ��}�!e�*�+�5U�$�Ӳeee�5d�IE��RW_J��1��F�`�y�_p؊U�o���T�o�I��S �-���� MM�>-�%��gQ&
^7  �6 N�Q�m�l���?���hdoFS��la����|m�&(����h�\$�'\!O~
��gąν_�<\kG�4�f˲ǣ8A�cc��~�G�\��֊YF���7�Ʉw4��΋���?���w+��r��;��=RXmI��ygP���n�PJ�uyttoM�/��[��Nw��z͸:<:.3�@�f'�� ,���\��?g��0݂�Knok� 0 ��(���D��(/�Bל""��G�0|o�S&�L��n H�x��6�]�]�D��K��O6��/	���d�bT���j�~���B�&�`dIP7�yID^������8��B"��)��|!�!�6�Z���E�����	?�y�ڹ����殮��3bOZ�x%�O'�܄�4dW����8��N�MMM&ו��2�,7�����׍��/�O�6�!�?{�U�Ӎ����13���������Q���D���PJ��:4jbi���N:�9��w�9��$Y5n$�{ʱ2�r @�4����g�zmx�[r���iA��y��fb+�
��)��[�Qr����c�o�j_Ix�ɐ�� ��t)���ߘ�� ���q�k���
X&b�V(�q<(xUQ��H+\�����\{Й�;+�󕦤����,���]��}�|иA~���
9���dJv��lbb�����j>5����d�mP����󌗉�|M%8�9[5U��������M�O�c��P������mh��  ����w��TѺ�������7�/���3Õdߩ)�X3��\K������+���S�h�g�H�������}v�=�:,���i�{Ӣ=��VewR����E�'�V����P��t��t�r�Ó�!��c�۝A�e����#S�- ���쉃z��kSR��īL��# &�a�&�I=����G��$�1YA�U��X�Z1	�R��y��JN��[���p�-�C�����Q
S濉w�D�٦�{.�C��o�q��P3Oyߴ�|����L�uF4����ޕdB�9:���b�8����"�%۵�����03{*?�vm�@�ę���2^s��D���p�LBs{�qZ�Գ��񍍍����[��|o�/�lw��M�5]_q���O�U�cjr]V�F_�x��2�SL���oZЛ9`�<$�BE�^�z�y��ʄ7�F�Z�'U�S\�*l���9�J��R�s��6ڒ0�����c�F"n=�"��;2����_��i$ҡl���k�-<���tAP����R���Iܽ
C?F"�9����A���snnn�?,b��%܀I��1N?@
���@z��E"d��ii���LPt��{��3V��>㓚�\��Y<��^�U q����.0�:���$��	���r�|�ݹZS8
�P�3c���_���Ȥc/{xxԮ��Uk��r����py6����U~�@2���]�ƌz�W:(,��TO6��sۻ�T�a��>�z�y< ULl���*�3��0\ɢ�����-��@"`�-�y`cRkp�1�Y�4la[ZeÜ�IhS���'_ښ�R�+t� h�S!n���#',f��߸�MGn��>Z�YY��k	�t(rd�q~]��A;\�=\�_��<�%��-`��KD��)s�Y}���8F������������;���?xˍ�O���j�C�R"����R߼�:�H���`��w�}�p�X��%�s�m~�h �h[U(aǳ���V�U8���L	?��$^��C�[�a�J�V�'*�~�͓��0b3��&Cr�m�ڐ=T#St?� v�^����#�0)YY�*D��ڀ=�?go7ra�Їԅ/p�����ek�ExH2hMڸ}���{�Y���R�d3o���OC�sG\>o8ס�Tt���6@)#
�j��"x:�pd�t�Y����V�L�J�!�O��}�Mf2m,��U�%:�II�8�7m��Њ
������[{{��=CjU�Ȃ��e>��t��j�y�{������_ԢG�5yZ��жR��IIA@dTR�7 &;�9�Y�1�� �¸�o炤��������)�s�M_)�B��M�p_#2rq$����ȗ�f�_%�b���#�����dq����s�!�B�_A���&���-_v���;J����s�
��r�?��6E��?nA�|xf��U$5+���$��Z����W�o�B	��[,<b��ҙ#F_u��"dX�F�Lu�&L�UiSE�-���хF���V�li����7r���_4���B� N�����z��A�����W��a8u�-4�3��30M{ذQ%�b�J��p�"H1?0��9��r\��k-x��	S�yo��=E�}��_X���Mq�A�ia�ez��%+�/a.%m�W���({���0�[ܤnf���w�I�W����I�����f  v6�e��o-�I�S�g����^H�HBw�j�?)v�l޼G����$DN��7�}�p��K囬����sk��u�H�"�| ��?�|���U�PD"�ޤxi�ono��$a���N��E�	������C7�Xqi�.��0���>A3��y���B��_MNR?�WV=���{�F}�N���9�~"�+@���<}Dw�iz����܇
�9���>ZT�ԓ�8`I�~�d�8ڨ?���I��MMq��#X6�R��K�3+<(W�I<�a���#��o�!a��X�Jbŗ��h�ݚ�3�֨��6j��TZ�ӡ`v��eE�_I��N(��"yA@��*�}��G�h��~��E���D4"
`��m�FN�C�Fׂb��ֶs��ε��ʞ�.J^`WN���9M�+�eC�j޽< տ]"�i�:->Z�r�끪�����d��vs���5"""1�u1��ML{����.��K�c9M�Щ�EG��Jы��P=65��z��AAo�ϥ�D.����w�R�q�# �C��]�����V«o`���;�(�8w�
~b��K6�$(�%.ҧ�n8�,r�y�F����b�)oVX]�e��wO9��J[_K�|�U�u����Y8;0/E�X0�I� '���X���������V�g;_�^"!����c����E��[�~~��֡�m��M㘦���tY�|z?9P,ֱ�tK�="2��K�0Ƞ���U=��1+�9^9�w)q����p!�����VhP���%�B�r�Ҡ���P�vT{ �P"/����o^���R�l�ɮ��:[������t�Ö�'(ׯuE([C��'�Sь±��*���Fq���X�ߝV�P����N���\I���MJ�G�݋MIs�q�L�Z�+Ѫ�Y���?��Ȅ�]D,"��M��[����Ƞ��� ����Ѷ���#��:�s������z�?V!�����FA�(l��u"]�z]���id�:��BC�\~/7�J|V-Њ�1+��p���������Ty����|��Ifb����4����X� � ����Ŝis����`Ͻ�-N�T�\V��l���~�lH��b�$5�����B�0~�L��+x���>��|�	hc����ٿ�0�����?L]w �o�?H�"e�
e���������u�Z$��"��ޛ�	�{�co�w?F������<�}_���>�纟�y�������B N ��0?�2A��:�A[j2I)E��c��!	y�䅬OJ�r݅�9+#eA����x�bI�[�ۇZE��V]\L�����!y��ȱ����/�0Cq�n��ϿZa��sS�V���i� ��(�����D�Z���T�I2H������J���ӊԩ�7�XZEj�O�N���%9�"�i(>�Y�>�&}w�Vc��c���ʫ����G��lm=qq)I=����F�J�X�?�7
�Zpl�U�����8?�U_�{W��'�D� ��.�h�4�A��[rW�v�"�<��R�55池��ۂ9��`z76uy������pb��Q�?������f=ͥ�t��Fp2U�E�������ra�ΠW5�z�����cV���W���"n��%I�A�G��-�N۾���%���|��g���ĒB���\���u�P��l.�Vc$=�
�3�� 2尨H��d�u���Vdi�w��9^�!����p�nYW��g�a�c�E��E����N�o�y���>6����aOq�Q�U���S�p�����R�K�&Z���K�N��rw��ݛ�6�/��ι�}@�r wKd�SU�����	�ˡs�{s�%���V����\����}��⢓0�mq�� �;��4bill�3*�%��/�];]d̹�z��_�6��;h���ϱF�����kV��:l��:�^b���1�'m��INX��3;>��}���'���N�f,(�P�������ߠ��|���oJ���k��e#N�.�����#�����>p�����F�)���:Ar���:�B7QL���g���)@%���N*~�����#f�����Z�&���Z�����S!EMi_���V:��#��Ag�*��l�*m�Qz:��Rݲ��?ǀ��Q�>��KE;��ay�S����_�����W��R��iR�}�?2�o,)��xa��Q~�������+z���,��	��U����f_<ߝ��J]��+X�.i���BEĤi��<�d�ykng�;�2��ZGV8A?ft���p/5��oo��ǲ�U'������s��q�n%�wwu�v�׌C�)��wZ�1��H��E1Sc˿L���"G�1,.,����mF�?�{Z\X0�X3��9\�p�W7a�Լ@/Ƕ��M'��.�|ys<��<F:�>sx�$���0��W��l�1��|Q��#���0�$m����u�X�ګ�)K���-���M�>�Yl��"�����m49{9�^�s��-�r�t��s���R�o_<ӊ��D���a�G����Z��>��S�����$��%a�����K�
4�Y ��~���hG���=� �Dٳ=�'����7n܉e�*-5�{c��I1���|����)ނw��5u�Eh�-/{u���� 3��{��9�H]/��Hmm����Oyo|0�ߤx/u|�rxq���UQX�h@c��������[m�:�_TI�>����l���H�s9V��0J��vN��J��3��O�U�Dd�]�u>��c� �Cq��b�{y�����+R@�8�oY�`&�٫� <��b ;�:�U���=�'�k�}��`ɱF�PS/2/�ݺ�<�����aX:���Q��vdU��z��p�CܡG�ŝ?sx��㎖��Mu�Ń�� ���(����z+7_����(��v5[[�����3��K�Ci���1�_XAO�R�������j�^�[��8�!i#h�*��A͒:[�����������\�e�ɷ�̈́�u��|�߽#�d=Y~��Q��q�m�퍌 :d�����&�ci��lb7�U��V�A���%l�$�-�����q����z|���:6��y�<�H�'C���m�l��=d�ª�D�c��KQ�����4r,m��	Y�@�t"+���h�2�����.�0:����~~8-�^�`�Q7�'z�_srڱ.>h�#X��"m�q�;ֲ~K�Z��t�,� �ǹ&2,�����\=�U����L���i����R�.����ݴs,�2��K�lw�˕ɽwܫK�71�&����n�O��$��	��)?�*�L4��HU�a@�P�Ő�8�u����?�}o���[���I4FA��
���z���d�uCܼ���H,�hr_#�����m��bF�o֓}i+7��st0�;��kk%&׳�C��х��J׊� #��S�{�[�=�RI:)����ʊ��5�FS�\�e����q縀�{`���>�Y��U��vS���){izs�,[��~����Um.o���~>;�T[���۷ɉ��w��ߗIWN,�����h��9�Gb���O�E]x翕�(݉H6K��'w�wF�k�����.E�|�0t޳?���>v:�'�f��?0j��o��7��f�z>�=ꖧ bk<09����AN�x|�&,���Nd����'�����<��K���-�4��)�	�W�g��'آ���쿲/�͞O����c���\J��9��B�Ky_1����H�����������:��@� �l�<Z���P�@��qA�`T��"���Ԍ�dVUv����P��Uzn�9�UzN��ÿ��\E�0�v9��D.�,
����Ӡֻx�w|ܠpHG<1]���8l�35s���x��������h2�O6e3�خW�p��'|�{��tll�k��B�w�7���[3�w:K�u,p��|������>TV&�;�����:w��j��Zwi�)�*x�X�\x~8L+E֐���MP
֜����ݫ�\=<�������?��A~���@o}}�F�G��(���D���
R�\���9�+֞p�+i�T!C��I�N�<U-]ɫxM�+������i	6y����Z�N���:��G���_�:¥W.�V����:Q{��1�@%w��%ӾC��o�|[x�0U�p��]�P#���l�bDDD[�ws��X�\*�*P���FFFzg��
�j�x�zOq�b/8|]������t�.�CK�b�VI<�&��0�G���<0_�T��έOn}�����B���V��3��EΔ/x�b����bxr����ҿ�<�ĒȮ������Ci��l�˰'w�B)�GG��]��������[�3w��wv�k�R��'�lj �yf�K��dp=�W
~n��ZhYCS�*E2�j��C��M7Й�M|]ǀ��WB\�7"J���}�)�]VJ�ӣo�xq@�G�d��`}�����N���I���iV`�ul�K�r�޶׺ �j�vi��o�ָ�o���2^|����[ZE��������3���Z���� ��0��r�"��LR�<�	�^u��ષpj�-Y���lfث�� �9��ڎ��`��>�ۮ��ԶuU��^�����$��:9�U�>t��ڏVn��%���Q^w��#��!.�(��z���	%�(f��ş�v�g6�P��x%T��v���kZX�}+�P��M�NP��M[b���'�(Ӿ%*�ϿJDd��ibec��]#���Tg8���n~�=�v\���x�{@�W����
��o A�3�(�_��g�ݫ�B���LbJd|�-��vt��距�<��xb]~|����e�����\���TogѦ3��Ȇ�x�Ig����dC��ً����姃�>�6��Jk2��� H�և?��9��.o��]C���"�鿭؄x��*�7\i�w^R��AG+�p>U!��̱������D�!���X^�P���._�?�2��V�-x�%2;��5}������ݓ��5���b�E+�E���hb�Ϛ^NKKВ���f\0}��6�g��2:��2)_ZMu�5�� �)�QG(A�ŧ�(k��P��H
���o)�*�Q'�����U?���������|�׆v����CX-�
<ݎ�^��3{S<:�R��ȳW]s�U�u�5U�^���=���ݜJ��3$q{ 7�*�,,�ο���&�7����<��Yu[��gG��2\��~�vU����Y��ӻ_ϳ����(������+%�G�[����e�fj�\�{i�+�E����{��wm�����~jjj3=��pq3�_E^����M�G�>ۢ` jW���U��Z�sasw� �u�lP��B���	�RW�;��΀����`�:	�����M�3�X)R��%�	$�Q}4�e�_�-�*ɫ��,f��w?���ԋ99�^�.���b�	`�Kߦ�B�Q?ֽOI�u�ڿT5s#|���}�{�O��G	`�v�: ���;y&ѶU�xcF����vwJj�]+t�� � l��v��hy���Q M�<j���*
q�]��F�Ѹ�,���=���WVV�:�˟���Dp�ͥZm�8P��5>ma����>3�A���#S�����^��h��D-��2�<0�C�^a��C�{�JF��`P��X�M�:)�&!�D��pM�q��_kk�Q̰˕�!K��˜��m�x|t@��'��(�$^�ځu��ۇ��Ź-1�����1U+�$�!�����6lP��g�l.�=vY��}�k2ds�=�حX�J�{��L�ׇ%>�
��>�BoSnpͶ���)1"���YT��<$J#�z��bуy��px�s�j`1Dm(U3.��rP�"��ݔ�nj#G�aI���e���/�c���z&C��C_҆
�-uL@ُ��\{K�~:|�C��-�X�N�S��˓�ޏm]V:�9l�=#OAI����+
���谪�����x��&�D\��ѭ,���V�a���C�Zk3 ���r���s�xǖ*XF%r&Dʎ��S��@r߇>�[���	<g|�]���r�A�QB�k&ѷ������WRM޽P�w��=��}w����>mGk#�k|�}��S:��؋u(�T���;���P�f	N
����orM]���Cx4وE�Wk�7l�1�yz��~��p5|i)�E�O\�CiX�OO������#�,#ܓm�U��I��A��,�? n�^+[Ά%�����,�����($1ٶqП ';{�z�(g4��,�Y���F���"mA�RHnF��񍍍2PB��+�xG-��㞈P�@�>L��P�:Q��I�7�_����W�,��s��ӍԶ>פ��'��<���iޑ��ɘr���lk�bֹ�f�9uy�kS�{���xMM_v{��ѝxt�kH�m�*�o�����p��?��2�lŐ��9���bKw�Wd�~Q�-r�x7{w[�n"�����\��vY��5{�Cȑ#�����~�_豰��1�h�@[�%����'�ƍ�^%���5T�Γ~��Y���E)�T�G��qJ����8�\)���'��d%<��dO�Z��ѡ�hh��������_���
?�8� �/M�&���23��*=ѻ|�~	�R	}~�άC�����{�6��p��s��U_��� ,�8��	 �,m�[XنN� C�xJ%�x�cϤC�xarR
8D��?��YZY4	���-�]�BYl-���k�$^<~:�M/�0�5�PDإ��e"t��s�Pz��S��&\��@���~�WYIC�̂�a�]eP3���?��{7�<Ѻ����). �>�#���+A65|ɜ�
L�[���7��Ɨ��3s�|�ʼ"Bl�X��:��Ӆ��,�A������������oҾ�UX15�H�"��uOO&���J󤨴�*3���و_U�Ề��� .����=�6�@-�Jш{�&��R��|ؔxД@ {�ǒg�#�9j3.���p;|IP���R�eS�+��p�4`���{�����0IC�V�N�D���H�>(�����iR*�9,��n����H8Ȓzp��n8��$��[�Y"�/^y?h��)�D����k$(7҇����$`�W=f�͎�k�x;���NΠ(t�3�Ƞ���;�8f�{3Q�������_�<��NW��zU1,w2C�f��������swM���~NX�?ܔ� �u���؎�\;Z]�f� Un9+;{L[�@P�"�P�m ��G�|ŗ�ķ��Fp2k�3]ݑ��-�ƂvqL�����n}6|�ݚ���~��IJ
��DӮMY��N��ϟF<7[��8 �j^m��:��n�ƌ�ݾ�bm�h&H�����W�b��d���1t5��
�u���._I�Y|4��A(vC"����ȥ.8�q|��[�HӐϾ26������Q��\��th�2^ޛ�>����W]{r�2�=u�Tv?'<��XJ4���`~�H`
�����<$�`�,�iJW�W���b��3*?D\ځ>{Se\1����� x��G �gq�'W}S8Kx�哙�4��&$q�����<��J���a@�cl �	0��8�������W zEQ��Hu*%x�fs����VJ8��r�9�;�S�,שO��7��o�#�4 �cO:{�^a!��r�KF�m1�?1�5y*|(0Z����9��n���.*��r�̠�A������:���qT	)�'�<����0K g+�s�p�|��3���`dPE����i�.���(١J�u�1	�:`jf�hQY�u %@�	�V�y��r���}� �m�B�abr�9���K���Wj�)�����*^b֢X���W�6U�,����
��"�=�T��m�!�<�KI� 5 ��98n]�)}T���d�W�2^�KxA�|ff��	d��X����bdz;��T�����k�~U��b83��F����V��)�]$#{"�QE�)�����h��'�\iDف�i�:@`�T]�u͇b�{�˰�������{{MLR�7#�A'���m`d$�,ыpw�EƵ�p��fO���o�%�&�� \�\E���s!��bO�3eX��0�*�p��s2A.|�|u����I�G+,�!:!��R���D�D�t���v�\ms��RG�Ē��б��`1��	�o�h��w��g��v�
?Nb���@~C�	>h�3��җ����K���v��=`%�F�@������/����NáYy���^`9:��WhC9�*W���~AL��'+\$ Ё�>Y�9=$��㸪7�e�JK��>\t�:�6�/��p�7!_������<����s@A�$
Wr ��Q]��)��I����u�.�����@�����s
�o���_Ck⁍�х����ʿĢ����vkpW�W����V�߈v�<[9���_/��U�K�5)�q%̊|�Q�{��R��ng�7 G�Ұ�ڟ`;����d|��ĹuH�umT�y�Eؙ";V~��(?�^p���[�����R<����%������'c��C��s�=�K��~K붠���&�TU��~�X)v2`>�T�Ar�6�Ü��>k�����Ү���]�ȓ1;L!W��yزǾtF�O���V$��5���	��Ȩ(J��J�1��Owܫ�={��:�\9������8�k�Ve��h�rG3s���N}������0�jm43�oT&�A��Bo���r�Z8���^۽=�U���G��߿}[*�.����8�ZR+��=�@5��x�z#� 	\����M���b����L٫H��oJ��Ûz������A_�J�R��0\��S9q���tzg1W�~��Suri�o!8�ψ	`2R�$.^��^3���XQ��Sݏ��69'�ݓvE�7f1��4�_ݪ1�xȯ���>pU�=IXa'Ш�z�0���5��`T� �^L���!ШDԫLp@nQKW���(����(��a]U�দV�v
�П�Ӏ�C�˟O��}��Jx@C/)T���Z�����Uw�Z��0��É�� �؃��[j�%�ԟ��l��&�¸ve[L�g�c�_�prq�c[�K&���989�B��j�@�����t	߅���}�~��1G�N@�g� �gz������[�h��!��x!VN|�m����ޔ�u��hPTgT=҄B>��Ʃ��8	AA�����&���w5�H2ivv�zH1���M���555U ���pm���9��W�������S1�	q�`��ga��l��,�uw��
8�@��d6dh�ki?[�h����f�9GM2g�SF#�^�r�}FF��Q���E�_\x454Ƣ	��A����Uq����,���H���쀸����I���,�z���Zw69nv���
�9DY�זA�3�ڟ���a|��X��Ӝ�@���?��S�Cz��|���4z�i�(<����WݍVe����p��Bn\:��m��p7�2L��Te��f.���5j��i�$�h�u�I�ߠ=�������9e�!ڼ���X
k�p"��쏬�W�I0ŨnL���hd�)�?����ax��юL����z��:nB����o<�l��Ms��j57�(�0ɒ^ʅG=f���R�]]]�S�p%P�*�W_��^c�h��<aUfUz���$�� ���<�W��|q��yN�eQPPD���:��YD�U@`��	� v)�8&�N�$E�h���~eZ#y�&�qos��{����2J�t�*}[�7���3O��,�]���g/�	e?彉��)G-Zǈn��
�Ņ���Wɬ��K ����qm�2Rͮk�����յ�r#�E�|1�!@{��@�U�$��ܱ�/�@Qr"�<���]+R��hx������
���Ӥ����4P�}N �4JNՎ���h����D���8q����l��Wн��剛��8�G�HIӕ�Ӟ�솲�CZ�~v�t�*^%҄��s�4���c3��l��K[�`����I�����afgLQ�ҍ����5l+p�����B%��V�4�V��F�4�q�6M�t�+��O�6Oy^Vu����H6Y�D��������9ˤt>�y���b�A�i����2��|ד��m�{��o��ȼ�F&-%�u�9���:y�����h�o�ø���G�$�[V�ҲR��!&�Sh�\P��Bֹ���pB��3m/?�b��j����v�T�t��E��Dt}��5�7��i��}'�y�J����G��p<�'�<����QL�i�cn#���������[��FF!L�	\�>snv"��=5J^�L���&-�.��d��	"BP\�J����X���={i�+�Gl���M��)x@��Fw\w�#��;�
�Ea��nޠ4�Mki[S;�����vGa��ۏ�.�N<W~��_��o�N��@
���,�Q�3أ[�{ȳ~�S/{m��K�b�A��r���N�)�-T���~��b���Ch^�;��;gyo\��祃�%�Q�#��'t����?�Ot���5��~�8b��,S>.���h�K���A�!�a�{��B�-����8�Q���-���K���u����a�vE*�9�8�69=T�YX�M��$���(�MT�K����⶚�/Q���k�ϒ3�Vmn�6L,����V ��G�}·|FtmZ��V�ڋ?����aS��l��3�ڟ���0����*_�_-�r������ae-{�@*�mj���َ;�6�`!�ޛ�w�9a�Z�
���5+��Kf����yh�~����x	�	�L�FI�l>tt�?u���#?�lv�>2@B5��X�d%������Ѕ/�4� ��ɺ�{��:�	dD�W����~�9l��Iz�\���RqS�݇%���Yc,?;<�G ~Ч�:7yU�?_: _b���cM�^���M�!}~�='4���9��o�U��3G�W�C��T$Da<G�˰�z�:E�<^䨬����K��'��#�.pE{$.%�m1	�6��K3x�i��{�$ܡ��)f�o����GzH0>���.��xm��p2f�"� %�ڑ��`�CI���w���˟�I{���1�J��aP�K��m�+LA���l�ڠ�:��}��Ԙ�����ɬ�V�7�r�d#_Q1�I��E���(~�91�AS�u���[����#L��A��-�%�f�������{�-,؜N+����[L�1v���O_���|/��W��.=�ڡ�#�m���@U���Fm�o�d�*��\�UV~�������،�j�n�?W�K����59E�/�6�tt�iQ�1���'��<��`-}���Kb#y&Y�k�b��oY|����#s�_�k�	iVI?u//�ne�4M�
h���SCp
�ĩ�Jl�0��j|'1� ��E��B����U��!��S�B$Z��&�v�w�a��i�.�Mpt�%M>�w��bW���Td �d#���Ϣ��mc�%�	$#G�go)��}��1hm����Ԟ������YvŽ�8M��6�RY�� ��9��&<WsK��d�Y8&|G��5脋���_�/���:Zr,�f�&���y|�$��1@�O��ɤ?	7�[v�i���]%��)�-=�})�U�_ޣ�on~�H%y�Q
��l���ʅ��&uM�����������wRq�bZM3�ts�����ł�[�(p�Kucec��O�+$fg,K.�)���,�b�7���Q��7��t*�ו�s.'��zj�9����s��|���_��r��h�G�E����=/���qN�P�*���!'��!KY=k.N�����>im�+������<q�̇��@7�O����b����@ ���-���FP��![Gk>2���G�+Qf���p;}����ڋ�z�_y\�37�e-��+/��A�)Ӣ�������~8��|�m�{@�츑���`��p��hEv����µ9�SP�6^ar��q�}t�C]^^�n���QLD��_W��^���:*ʬ��<'WO/.f�(�N���� ��ك˩�_��vFG?�2N���y~ �K��ؔV�7���x߶$W��b<W�����:Z�Z�ڔ�9����:�>���3- N�'�W�E�)@������*X -f,`*�����4I\1�%�F�*D�Z)޽+���/��7mJ�͙;��Ԯ����QߚHLk��2B�����jW-o���x���)ۆv|�9C�e"���D��[ 9��y�<r�>��y�FP���}~Ӛ�_���Y�M��/u�f"�ڮ��	�����"MR�����t�D�SS�! \���N���h<q���n8sd.��(��Q�M��g1)_���]��r��!�\�
�]h����h����+�usKK��!��������Q����v��ŭ�Y�b�L���@���%έ��v�X-_z	�ӥ����Zwnu3��+ �N_?*�2[��Bu\��Yo����(	;��B��q$@ hY���׻��(�5WY��`0ڱ�l���PD�x�v���N�{0�d,F����/����b5&���T�DFE�!a�)�"u�{��6�ux��!%2{vi�
i�����2E�t�Zo(w��j-����w��Ķ6�b�W��ԟ�60E64-�Tef��^���c-J'r�0�rz�� 슠 ����2�c��,�
ob��`����E�u��BXS�f(U⎏7��s�c�����Pfs`W�Oe��Z��	��FU؃��v˜*~bZ����'ح�j�f��&~�lP|�8��N��}:FϿ�ng4�I��#ڛ��b|��"������p�`Pl�̻��Am��H>En�����������+���4P�˻�TI�y����=����"���<���-����U�M�Jq�s���-΀��J!�(u��d��u65�;`�������b�
�j��Y�o+]ʮP���p!��R�ւ�_�E ��q��D�~��^�8I<`�{#5$7�LZ%�����Zڔ��/0s�OfUE�G]/H6B#�T�;��}��&�i��g�O#d����-�P��6����[��o@>�w����L�3����Z
�H�"UE3��yT1��q!;�����V�)�iKa� _�g[Bn�J*Ȳ�No�z�����i͇	N��uŌ�T0:��ίQ���}��e+��/ H_b00�y�µ᎖R!�����y�!i��ᜮ��]��&�f&��'|=�o;��[���v!Dd5 �ٖ̍����[�U���:6���"|�Y��W>�ׯ�9��u���---v��%`���|��6�y³:eXR��3���)����I�����z�R��'�	_ngy��S�"UȤ�<��1��g���R��Z�����l��Ͽ��I���^��C�Kbkn����\��1��G ��S�Vއ8�� �:��V�c�#H�F,��<�c�q;`+VY��_�ZĲ��n�SӏY��8����5%��9�E�Z|�͕�:\����/�׏G"
�`Bt�i�鍡o+�Ņ{�O��< �KC``����=�s�C�^��b�o��'��պU͉��?����lY��M�Wٝ��v7J7�"ϒ���y�q/4X���v�`�#Ho�Ǳ$���Q�D���4{r�Fʗ�S��%i�z(M���Nk����ё�����/FGA	%9H�� -��G J�+;='`�U�<�+���?Y��2`��x��}F��t��o�#�1�a��6X���2��}|�99�B���᪼�r�.�e�*7�ׂ,��n�՛�����Č���;Mz��Jk�h����_t"k�<�+�
�[�8��o�HWjƮ���֟�����_#��s��ksD� \SG�>��������e;��<��@�8��8�<#^�Q��M��G�V��I����ނ'��5������v�'{�����|�/�[Q�����������Yv�̞={@@�y�)HT�c�J�� )��L"��\���x�IM>��������6�o��o������L��:؎o�?�M�@�y�B�����d�cH��_Ǘq�����1_�pZ�
`���w�>���;J��7�Ҭ�2��������A�����S-|B�/yb[?�<m�U��Y��'�r��1��?{_���m��Ό�]��e�.��4�GSrx'���'�v�x%�mËN ���?~2�5�������X��y�!*�٣���b[M��ｿH$h�%�m~��?�J|���k��yNr	�Q�����>BS?�ÂǰG��T��g�~Z;(��A��:��B�c�V��uID��W��yp�yO���ڦ�4�1��W����խJ�抔?�	(E��L�g<sVP)�D��S�r;�ؾe�����g�5�Y�V�9�egGQ�>5z�Ay��HT�QW�j��<$�E���"5?=;p��ݔ�"��%���\J/�����_�h?Bs����
M�Xoſ4�ѝ�Ӝ��ڪ9J+����_�jg..砬�~gi����<O�����x�������X�\�
j6�V������,�K�9=�Y)ѽ���W .3���RV�s�41�w�1�0E�x�?������t�y`�h�t%{�������~��~P!o(������Y�ҜPR� ]������_I�X�q��Q@2'������?�2���R�P�}�c���NN�ْs8���ׯ.,������v�ќ7�N2��M?@�?���&H	�,��٠�*X.��U�	���		��\��&�����,��(�Z��m
��f��P�d��{avRC>}�劋��`�;�o��%@�@�=�v�=�_?��k����E31���%��/��J7Pm���5��2rY��|!H�����kU?=��u�gfLүa�\EC:́�d��*i7-�Q�_��=+j�Qj�*+�e�M����M��	�A��y�g�k��@�k��~ D�(K��KL'�EX�"�;#��QC+��q���c�J z��}���w|����. *��U�?�S+���m�� �a���� ��,��=�� i�έ75睮�C��[��/Q���LOO���h��:��b��	���c�� 5�g�5�5��g��]�淐G�)�gg>]f��e�)8��1�O��PnL��:�l���5<����]���l�G��=��pe�ha��~��<��`$
��F��c�6�?��@�#@��5�Qg^��B���7����9�Gp�q���߭#i*I��͜W��4K}�Ӭ�e�#jw�L�����s?
��$b�#bWڭ��l�l�����Ȣ��|$�r`�2ͿBЭʚ]J,�Y�zM3ѿ?ބ�D.�&��wi���h�.o�/v��+;ލ(�N���X��R�t՚�ݨS�Y紜�������E�[U]�>��(]zn������ Hy=����=�(��Km@�)~����B  ��M������hdd�TFz�� }o2
���w Nbn�T�2-���mC����;rHJ�����+%�	�2}��<i�`��C�t�7��\O������+���d;�?�N@��	%vӿ?�l A�i���^Te���wә}���^�{E��$q߳$<���A�'��n����� ����|kо�J>z�ݛ����V�$�A�҇�ӹ�:-k��<�� ����힍S�;o��7})M�J��5�v��'�k���4���' |Ŷ����wV���e����&J9�z:W���3|B!C��%W�����c~!��x����LD�8ڀ��H�B} y�Z�~S�L���T��� =-Aa{
|��M�ԕ���B���~�Y2�H��O�� ��4��a O��S�v+E�i!�����Oy�����{�����l��*%�K%�Hs2���;jÇ#z��3�5}9� =�S����Ԙq�wB��e6����b
�`�?�ޘO	m�3B�1�@�+��rr�W�;#1�8�:H	W%9V+֪]'�@�o�mЊ����e�� t�+���9�NɎt�ջ\29��v��#�r���3�vÚB�c�#(���>:����yU� �(�VVVY��(�S�D-�ۆ� ��G �e�;�(PQ�hS�f��K>P[ŕzaS���%]3�L�?�%�b3j`�X	G[���0�w #n{^�_B�s�� �x�aWJ��c6���.�C��v(�(+L�qx�h�đk%�v�|�
�A"�k8���ޱ�oV%ܔͳ�ې�Aw��(deg7B�\���ux
^����i&50-.@�쮌��JM�
'x�n�򾯡�|�v�,Y�6����3�Z2����:����FA��H@W�8i��a&u��^xjJ	4��ehV3R`��&�{V�فʞS�2�
e��E��%Y^̩�d[�-��%u�ē	�}}���&�t�y#p5������`=6E��$���x��	b�O���6�{�=��M<��ˏ�a���_���6��"��
�BB�'�j�*��i��cD��_T$��U��c&��`�*�Fo�7�Y��|3MN'Y��������P����prys�	�8��Խ�QP�ޯ�rs��yقz��oP����G�1��yݶ$����M�J��+~�������#1~�KS��/�98RC�6�;� �=w�TY|'���H8>-�]��v���RЈ��4�hQ�%���]�s7z�����cy�`b�i�p,]�pA����l�D�aVN2��`�M)�>n����;,ymF�\�,��10�@W1��zJ-q�)���ݙ�߬�h�Av4����Eԃ�o�!����SL�\��ls��UCο��l_^�~�l�8؆W�}���� T�y���u�)�`���6?<�)������ �ٻ=��3;�7@�����eu��Ln�'qOz�DC��+��+>w��E�,>���O�*L�{wz��P@�P<��"�&R[��q���uAB/�:!W���wc��6[�ڐ�XT���֌��$����/C�]�v���hhcA�G�)H)V)��kщ?$�"T�H�#�����3\>�+;�����^�-��7V{aTe*WL�n�ڃ^��_&ڲ���t�&� 9!�3W�zo
�����/��'yȘ�1�Ml_ll,?�����7�ӊ������i���f��~G�/���j��JC ��N�F���B7�c�E�E9^���O�JT*����n*��؜Au2���e֢aɏQ�^�jv�z.@��)@E���NUG�C�HgN��ʈ�3�3�}7�[����A�Y��{|��̍Y?~��W��	��}G �~�J֖���W�<U�4�8AR���� �/ ��Z��t�͈?֚c��K��2)��~N�r�pQQ��+�^^s��_�dK���6竏���iNֽP��ۆ!M�4�d�5�]t���B+b��������۫i/LHi��Q�{���ǡ$��U�Q�)��C��c��ߦ�b���G���9���㍔��-}2i���,��9�#�n�(cM�=�A�\bkq�	�[��)vu��b�=GB]�����>\3���'�Q�!��)k70'���(ȹtg��bpd�'�j���v�V�M��䅵;�rw7�g+"c}��N.�B^&�%L�\]IFKE��OL�um�Յ��4�H��?G�Z�c+�ut���[�*�u{�~sۚ����_���t&>���kj�#yS��>}.V�}�
��V�Ì�u�eA��V��e��'��|�/68$�^�R��d�oꯉ�}�iW�C�-w=�ܪd_c��kf	n��3w���VM�sz:�����-�X�W�Љ|_qMs��_?pU���	O�_����rGv�jQ��z�� Q��xu�k��5����W+��W��y��/ζ�Sgeee��*���|�J	���6]:����5ve���E���p/~����KGKK�]���@��3U�/_��
��|��Y��o=�ٝx�|n�p�R�ѧD��݃¶���	4�MW;l�col�!{@qqq�����JT�Z<]�ݟlv�J�4��0�ӊ&)%E�ű�h���x�X����S��x�l�/О�6�C�X;x\Kp��<�zE>���Cb!�m������ !��o	�M�:�'�~�����������M�>}
B�;B���OG��o�{��ӵ��d�˰}�O�z aF�豮��%I�k|���^H�����!d�!T�ԮE�g���z�����Ż$t��h��њ(!14<��s��"��R�Q%�ߝm2_��p��w�ށ���<�`No&w�����)|�wX�q����$b��߭�1k}i@���hvj�kË����X��yLVS�#��$��W��Т{jġ=��׏��K���@��,v�UC�jj"�/�H!G��!i)7g[���&�HK�Ĵ=<<���]�`	��Xt��G�T6����m1�;�z,���v!��%_���k�Y�Nݥ�T�����3-)l�d��B�VW�kdi�;99A����V�W= "i]t�|��g��
%⪼�� 'C�j����/�f��o�10��w��h
���J���3p+�����+�K�#"�R卺�Ɂ)O�[V��O
���TS�ᆃ���L|3�����2������Z`1#�(@�Qv�+�sg�N�u��ٺ�����UA$#��RU�ɾU��Ew�>��&��C�h&�
Ʒs�����Yd;]��˃�h#BJQQq�Mן��ُgyF�������n@=��w�\��ǩ����O7$�;/@�*R��9���c�M{�$� �&�vp@^�d��ONNf���ԟ����0=@�m/��$BSиM�딦*����n�@ۣ�k�r�t9�%95�ֿ�2�#�����x�~东�l�7iI~�ؑ����s��I�����ј�X���Q����f����˧�_D\l� ���?�'��RXTE4��R˕����Ȳ_FMM�=Z��?�gj4|�o`����$tKIl���H�م?qT SH�<W�	 ��URd@��e�Q80�]�{�R��Z�.��b��S���C��] 5e��������w�r*e988������*��E1�e@2
��
*�s�DE@� A�E$I�X�JQ� X( YA$�R	*I$IF����t�s��9��ޟs�{�j��&3�����1�Z�/�h�S����;ݥ�%iHt�����Ne��G W�!WD71[C�iU55 ���R�֦^��Y�{͌���{BL�;�|���x�n��76�
�u�x�]^r����M�m�/�'���]�-8h��|��(�7�	Pd��5��O��qAB}�O�C2J:�"5x��A��`pS���ն�����
p�}d��hN�l���ȕ�u�_���Uf���v�up��ŎBo��))���C���"P��G���a��P����N�ԕ�����]�/ $���Pf�~�Ǉ�jj�?vm�����{9)�������p�R��/���6
�±�h���|��p l[:�����(Yߨĳ�7��g�����ff�,��i�	�o�wE{M7�J1�����Vq��Jiizn���{_^\z��h���,�0��5�*�NF�����n*q�`�Y!�+����'J·<��yݽ{�|�5�gֹ@�� �h��.Nj��-:�iu	�4��ÇU*�K=P��7�XI�'J"��7:��7��q��@I@�b�#Q��b̞����,���o\ؘnF���a����; yV��ǡ��	�g^\%����?��m�����F�ۛ[���w�!��D�%���O4��C)+((׻��i@� NMj]�K[y�N0{X��Ā��l���6L����l$�h���!�jOq�B���_���a��ڐz����=�	�k	
�Apz<r)�Z�vOy{��������P\T!�̶�����}���7�RJ9tu.���Dy�6A���t�p�N���ӟ��:z����������uTJ�4��2Z�/�N��%]Ȉ�X/yɩ��?F�q�raP,� ��(����]^�}�nb�7k��i>?~�Bsf�ʡ�rʻ
�֬.��͓࡝��,vd���0(���֬a>�t�<	rQ}����b-Nr�Z��9u�9����6�B�t/�!���<��� `�{�#]����]D�L���Ij*�Tu��/��t�y�g�B%����M6�^���* �;��L�����]���ڔb� gjC����u�&�nnn+�K�ښ먯�펽�utt��g��d��6�z�< 8��}	�hW+�2_��Ն��������v��}K��|��`��"��u�LϷd�����S��8
�B�;_U+����P8oC��p�?MKK�g�tV��<���ƫȗ��s�:�Jr<a*����{l�եw��D{�in3_;F��%��mv��j+:-t藽��Oq�o�P���u�ߠT\IP�ם{Iq���~­�3�z��nQ.jβ1h�uR>��{�~���	h����?���x�p	ڬ��mg֧��(�(������4�Tܞp��՗�{��:�{LX�Lo��������EU�><�s|ݷ����/G;I�ػv2�y��U�꺪��0�X7��ʚ��� �~��.��z���
��S
"���N����/*���V��ԟ#�|}g =�v��[h��l�N��3_{����(�TVr�0J��%��� ���|7�>͑�m �bߟ=f	�-:bj�k&�	

B��:٥gN�����������ݭm����`�_܂P7\��AGL���]]t�z�g�9��	,��(��<v�~,��jӗ�"}[[�� 9��赆���~�a�K6C���kٚ�H���A��4Y)�I��j�N��N�B4!ޝ2LIL�<�bl�\�R�P�N�������l��.hWp����Y�Ke�.�ԉg'��W�Q�, G]]B�y %o���Q� 1�.�\�+S�v���P*�C,��1�� Ud��)�n��9�L�L�2�?!.�Ƨ����;k]��O��$m�&3
v�T�i� c�[|}pN�%�����ggg��:Z�[��<�n�"z�H$�^X��er`�K�=�+�9�S�X�����%)�	ӋS{�������zܑ��<�2�� ���#�op�411A�+�G�窕Q�L�ϡA��M���90oA�������؉��X�QgRUJ�[t��܏FQd�.&&��5�;@F�?����������~�3���!UO�J�Em���$�䬔�^�a��;���٢��0�$��yg���~TYϏ����wBѮ9ˇF�o߾y0
�G�����	��p	 K4������߫>����(�/vbA�5]m��p~MCd�ʕ�[v�n���ă�`9�;>A)I��^,p�������9)%�(��o\�ˆ��7(��-\|(6�ڡ���Hɗ��15i��@�b_�/�]�L��1ӓ�0��~~����T��h��"�P�������*�ċ��VS��N>�S�c��w�b�QJ�ph��@ݾ�0p[��&����̇�F����/�όw�?��#C@u�[��{'�e�bR�)�-a�"�O��?��z�}k�CCf�~<��,��FH4�Ywȝ�؁36 ��}ū����]��n�?݉���(q�/���N�}��sx�]�9�������KÝ�.�~��k� �]s� �Q�0��E"����)1qq��欗-ٙ�n}���<���~|��>=�rs~��Q�f��^m�366��ڢ�:Z4=h���ޟJ����ڲ-��	`,亮��h���;MaKs]��mTV�(�]UQ�:/�ܦZz�u�H��8 ������W�v�(!p�ݻw��س���nq�V���@E�{J���4��	7�^>�%(%F����-���o�������xqq1�f⿽����|Z"]���'R<v#$ ���a@��a�@��H�)���'�ԙ�~��;��Hî�~.��FI�
=eA��g���F{�I���������2I�\��⑰�nY�0��S����=K��!����;���_N�8���+f�]�ho�vA /?8]Hq��y�Y�'��6g�@�'�/t�)J��l�~S%�tDT$�l��$����˖��b;F \�[^�07�2����u��s��},&xk�N�?;?E��Ժp�iz� ė�ci���$�<��Z[�iU��]�v��O�갧��C~��"��b�ڊHii�֎��ٳ^��[Z�RAA�oOn�|��N)ccc� ��a���}_��,����֦����k�P���l}r	�D�_�h���S"���fH{*� +*)�(++���馶�:���S!��pG�J42�����ɨ�>����#��"'	@lA07�4z>�B���0���ͮ]?jʋ���?�M����S����h'��+>�_M5Y	O�sjjt��U��.dX��
EO���v*I�&�H-.{���n�0A�Pq�������ʵO6�d�n���.�X�Ag��r�4�N���|�ɴ6x�{�c��f#�Y����I�ZI����ж:��|�;���^D�oș���u��6&��7��GBhE��a��ND����Fl��c��X.��?��:��_x}��0��_vTJ/�B���?
�Wd��ty4'!9yH,/�Q__�;������1��8q��?	�E�rt۠��+�.���Ru!`�Ƒ��ne=�=۶m�\Z��k��]7��8K1Kq]�b�/�E�C?&��#)��)��W��	)��`�����{�4��0Q��![dِz��U��R�����A�)�.F�qU��܉f���6�Ag+DZ�h,:����VԺ8L6�����_�n
	-�G�쵒cx����\gz��/�b�dz�p���0�oW�&���!,�<�I�12�O�B=���I9�/���SYC��m����&`X��J�>ϥ�9��ո,�ڨ�Ol�(�Ӄ���{R��7����8��kmà��68r,���Q���i��\��{0�:��䯓�N�:��䯓�N�:����ѓ�{��6��ݺ4��5��ţ�����t��c���������U�?w����͜�k�^��
����y�ê���_��o�o�p��N�[��V�~�����Ͻ����E���_	�%�����KJJJ�Vɭ�����X����(����N����&��������c�S�Ɩ�TTjW��ڸ�������I�N��&�n11�S>�md�uq���V�'M�V�'"���4uf �֟�YU3�u��~�����=�𵙡y?��>Ӯ���8��a��$մ��.�W�B��<�]\0�7��QO5j��knnn�.��Mz�`�}���ƟW�)k�H���&¼:�/T�:�pqq�V�2��l��ѝQ�UkP\�~]����8��:���TƂet�X�O���ǻV'X��c�=���b�����Ɣ����ʿ��K�/����8b1Iq�2�i!����Aܽ����$''����E�s����p�]eSS�e�����):F������!y�W3��{z�'���Pp�E3�;Mn�֞�MV���jZ�FT��@�0��������K E˭�w�ۅ��K��E�+[w�ۺ��e�F��[�:�L���ެ���?J�_	�%��_	�%��_	�?!�q,��zX�veeҽ���xh�'Iifվ�ȴ�cV:�?��N��8>�ƭ����O���s�*��_l#�o~A�?����K�/����K��;�$�<�R���9B��<?��˺���{�2>*h�c�;q�С#��B�_����]�_'��u���_'����I��vJ��#�9}P�l��s�N�|�^���������C�ˊ:��;���x�./|Q�n���N�U+��>��5M�z��bk|q���d�5�|�r�!�耧�����3��e(<e����Q�M�چ�s�Tda����!�%�{�8�K�֜yk��a!KA6����y���{��pݓ�X�G��T�y�g��"��):���z�z,~�GXNz�^=>n��vk<~	�+������b�y�ؙ8�Pۜ�3d-?}�:\�c�J�=p_��$���&""�L�JL^8����JZ�����ԑT�_3��Sxn���n+��D�����%8��R�ނ���r�@�
8�"��󔽐�n�\B���k��QG�c��_-����t�*"2R>_8��y�8����l�D��3��r����)��Z@!��U�i����ИCX/��`]�\XT� �=nx�U�9�#Ұ���a�Ǯ�Os?Wk�2Mk����7�S�����Ĥ��`��8f���s5
�)������8�,��o�n�#�ʡ��)��A{��o��֒7����Hx�3 E��k�j�CDr���ԏx<]�����H:E���oOi|�P����j�t47:���* ZD�\��QL��'�s�G����}_0*T?��H�El�!�`���[G�絉��tqr:��Ĉ��rK7e١���Oc-X��߮��!;E�l� \�_@�*�~&��ؼ������y����������J1

W�j�&���1qV�&�Fq9s��YZ����! ���U���-�3����_NV��l� .��dl�	��C�����tOn��A�B�Cb���2����#�����(����1��j�����+zm�4�&��ﭳ����!�]+B�"��_JRO �+�ayO(x�I�qe�9��a� sH:8�ow���h�y���j���\Ľ����1q����p	8ڢtA�9�$g���Q��v����D��L	��$A�h9/b�Qe<R�_k��	���v��}mNN+�H>��#I�f�I��b�wY�an���'w�"]�����r����?���sZ��:ϓ#�c�CV`ĜP�EƲ�^sZ�c?��i/l1g@�2�@8�g�	1���r2�b�!/u�r���p�u;���l%XQG��V�`�O���
�Ӓp�_���H����(�M���<�7Hr!���T����ɍw��z�p�_�v��,��>���p�����]��Z��_�E��q�UQ���Q�d.�G.�R06[�& +ޮw���,h ļ�)f�M\�u�q�Ć7� 5����2�"�쟝���7������!��f���,���S|x18C.���^TP%�S��8���,�F���w�<r�>��n9��J�Һ�bǑ��U|�!RL/ɉ����?Kv�(��9gD�j#.����,��i69-������X:�����x�w�������3��d���Zةù��,��(�K�vb�
ƅ��Ew�B�w:)ƪ�S!��,�q~z/���[[li�
6��0�zF�e|�Yh��B�6X��	j_8�L/WUp��v��е
ӂ���R�/�a�C�� <����gh�'.Ml�_����cd�m׸�J���l.��Nx��{6��. !�q�0|^�7Y����_'�\����Ts N|j�;�g�*%b�F�r�Z�KG�
���:�����.�
fB�����뢀�O:)��B?��bH�:�zV�̂�ܿ�q2{aԃ�U����+t�[���L�UV۟���8ƿ�J�i(F������ �%��WYp��m����a\sz�Z���^h&_\0�OF�t�@{
��	V�lbG��N��r����&����>�[�8Ym����b�?�ܽ4^�oGvy� �P��, �w�A��B^~���귰������Vy��<[��A�8J�*QӜȃ�������&g�"Ռɇ�OY៑���wf��'��ħ��$��〒����C쾝�r��j�������	�V~Аm
뺩������L�h�`c~t��t�w�3�M��>��V��8��cϥ�J�&���"������s �L7`��r���9��BAz�����~���y_`�>���M�`�1�ǉ��=�g%ͼ�P/�%(y����6��6ui�+K? 8O��7.�h���D�ry�Q�M-�zvo�M�L�y?� �cIc�b7��Ә��;@o/,X��y���Xd�qb���6ֶÔ�O �<��<}��%�7�fi�-��`��ͅ)O7XؽUؠ��\A������`�����a���s�R=�%>⛯�'���|g��H�ЫM/4�K\���\��W�}�I��>9���֦�ʣ���6���w� ��љ����k,����*��p�aFP�M�g�x��6�]DPO|=� 4f�:ݦA��u3����#,8���&��Rk�!R�V����=b���rWS�sL���J����A$X��y)&��~��������O��`K��j&&�����;�S���F`����DԼ�6�q���r}p��+�{dd rY�0�j�J���αm�c���Im��l
���!�:�g��%�7N�����L|f�1��N��z�+`;���������TCқ�0�Zd跡z�k�q
y`���i�X}>I7䔥�o�'�kz�Đ;�pݥ��(h�5=,������G7��Ɔ�c��Y�ۗ|]Km�7�k임�@��#�+�u������áa�K����@�G���H��Øh�=M�!���U�]�e�O|m�N��#��q���:���]a�5�Bhk@�e��@T+{�eh@�)��;�h{��'HM�ml���h9*6�z����S&����!�#1	�v���
��	�ȸ@��a+	�w����i�҈�ݗ�m��'fx��>�A�YY������v⵨�*�w��0�D+�Zr	���6٢Q�C��M6!R6��d~d.N;Z���e��\�s�YμfW�qW
�\>�����.���� �?�u����,�CO�+��ǧ�!4nm��pn�5��n&��/�;P�΁l��p��d�h�6�"�J���W@�R}*oB�,ݔK(3�}`���{�bsV��c���(�}��'�[�Ÿ�}��OQόb��Ȳ�b��e���a�Ox����C�hހ=�	�&��.F�@C �a�=��xp����'ۇ�������δ�|��7�6���0Қ��d�>����)��Oq!��D��,��k�B���rH�z�6��F7QE���d�À�BP����o��.��pֱN/�G��<�H� sK,��F7C^P�	���A!-'�;�Z"��� ��l��Bl��]��˴R������e���K#r�5�̸�������3����i�Z%�.�ݼ�߄���(z�ly�~֟}OT9��.�ԯ��G�f�r�&�hhvS5q~��s��n�X����(��K;��B3"��VD-2���"6݊ޮ���Sn���� 0,a!���������\�M@��+]_>����0�?��u(I� '�%�e�6w6�;V&4�	��";�__��u�)���_i��P�j���|nf����n�g���^�h��.���t$`���7���A-XmgIo��|�`�Nm���Ǟ':j��]���_s���*+��Jn�Q_�t�K}V�{���<�)�+8<��f��@^��@�|6�ЬCF�r�]�
��j>��р��֢艭!1Ff]���Z�0�z�?�tJ.��;@.짉����O�]{kA��J:�g=�u�\���k@G6⊯_/i%%�+<���b�#�Sh�	��ݏ�����lA�3D����~�j���RP�VH�d�<�����I�%
L����w��}�n_n?ǂ�z���+��ep����Y�S��R-j�_ތ�� ����3g��W���SX�˚�C�B�*�4D�pV�8C��{�޽{�/M(r��Al�G�[�\��.>#]+$:u3�'.5h_�"5���Ėk��vC%:>�r��v�f���'�>C�B�nW1ҙ��E<�����mL��pt����%0��)Ȯ��_M�q,Ԕ�a߲/�{i`�V]~�~����ǘR�A�p�3eB�8hܤ V��1�
C�1��ZI��WZX�>�'!i�*�<�C$����cx��#�YO _�;Ԫ/��� �Mk��{���@�n9r�0	�?��Ğ:��n�S�2�5���KƅqN���N��f#r�gwȸ��l6������!.�g��2������ܰb�*8����E���2{˛mV����{��Q��6���O�f�;�3̗��D�|�l�������N�ޕс"�	մ��$��Su�������(�W�7�o|�}(�3X��Dmt�Nb�q'-J�+΋�͞�U�����2*?�9�,q!�"�i��J)=y�-�Wi�?�ITWX�6r/a��.:���k��
Gq��k�r�uM��?�B������y0�����@�-IP��W*�}*�ȹ��!o�/��{�¯�X�����M� �S��
u����"���R,�R��0�]��;6���2���5Z��jy�g��e�ol���n��ij�� 1\�N��CF�o��>#�֣���,d<Q��	�IN�Ѷ ��~[x�6��yiݯ���rd��ŵ`x�]����*�����؆&�"��:����,��9� ~�G��������S�T�D_R"��k�$�両�Q\~��e<�Ϥ@|�A>�	)�,��5��g2�~*�I���D�瞫���j�V���������>9ՍR��߰��%��ʎ���02�C�����Mُ��ߡ��ˢ��΁��wq��I-�n�d�Wa�69��	D����-K�����E��q��Ap�<����f�S��W?C��~���~*�< ��	�6����� r���*8#����=N�t�*g��a�N���A���e=l�}�y��CW �m��yn�]���UM�OQ*&9�ǿ�q��Cv7�}W��,c�I"
����X�h��e��ot�ّ=�u[_5�`�B�����V:T��!��D��"w
��� �tr?����--�B�����1��{����d*�=�dԸ���HZrG�:�m�BJTI�nҾe��KȺ/:W���'�;Lv� L:��_�����n�����l�^&xe&=g�&-N� ���G	Lx6���T������ƵB}��-[���"�����+��\J��"�l jd�uS�_�X�cu��d���A��d�c����fA�Da2���'�r�5���8�\f��{yXY���= Z�~Xy[�5Se�Ĥ��o�P�.7���~�lHe�b�i���c|�ktg�>zzŸ����V҆k�O�'���^-s�ƽX9�#�l�*�[����Υ��

fl��
�Ė�?�/�����=�#6�wkY5'4�Ҷ��%��5���:�鞁r�& �q499?�:M:�q��"jJb"��1��EF�J�r���|��ŀ��'1�<-�w��؜2q�iO�4K������c���w[�ǘ�C�V@:���9_"��Ecc״����bK��������[���z_]�͗�l7���<�{�� �w�ǌ't`�i�r1�ѳa�l'׊qI�s�MI-d��12�,�u�=Ed��ђi�͸pq��b�����<F�����g%ŵ��O��?�A�u���~2I���V�h���G�c�k����N&��:�X6���s��@��A�bF�����cn����!�H���'�D�g��`}ExF�����nKI�"�FFݴ�3D���3�:}0�b�z�)Q�j�֍���ñkC���^i�
�ǰ�A��2Ϝ-��]�Q{�r�Sd��iG���n��OC��^7D6�Z��5ӄ�}͊w����ry�K�T������;�xVJ}�ll��8�O\�L�w���A{�+�H{fjP�;�+�$?w���>j%&%�*Ӓ���%�u������f�5a�շm��@�H�xll̻`9I�t����U����k��M�'�u�o��!�do��[)�W̽ON�\�15=��B�U�f�3�#u�L�
�z>nQO�B�=�>��M`h�-�5����ѿ\R�}1*����W��~zE��ӥ����E��-��y��m�v���:������;Z3���?>nD��]#��
ȩ���&����,xz$q�K�gO�E�h/��>R��l��:9��4u�191���{��������i|�9;����M�p�Zq��n`�J��+�q���*�e�l�ciJKKc���,#X=�Ӳ�!p�����'��Ƚ[�S�J���-�M�/�#X0�z��3M���L�5���$�Ϛ=ֆ�|z<o4��D��F>�LIV}�NTd��ǉ�B��L��6�H���]��M���㉿r0�;�]�"77��="��T:76�FyMLL����z���=���0n�B,EKG�O1֦cx�삠�����qvn.��2�%������g5�J�E�ʑ��i?&�=�o�6p�
�J`�������B6�.���c�����BB�Y�sXM��w�Qr�&���	��/M|C��MУJ�UeG��MN��]~'<���b���."0y��z���\�i_ff>BF_d��켶��fnn�>Q?�s�p{>���� G4��+Z�CR`L�v�4(���.�c��kkk��O�'����!M��kzu�91���bbb�q�#��*������ V䬦����N�!.��7D\@���2��I�N.�8�9U�	q�����t��e��\� �llƗ!���[���ϟUUDFՒ����7�r�1���{�����?T8�l�ZPw����Y8/:��n����ߡ�����&FF�ꞕ������ �= ,�&���%�A�˱�x㨘�8�|�E�$S�P�M}c��=����\�!��v&ϊ�����+'�^�\�¥�O��и1�+d�Ut�<���׸�Є�_м�2�^�(ڟ���-@�K~�5 �FH<����3����-��0���CLE��9}�\T��S�h�B����|BBB�bbD*&��(7��f������]7޴���Lk ��w���@���Ї�� K%��,����I4���Fsv�
;���N{ǯoo�u寨IܐX�~�}[fN�6WAP[s�D��Pi8z#�9'n_�o�~{��s���N��!�����RKG���@כ��e����>��K#6�4�ie�$����`_�'2y��/���^�y;{���͛7�a�;W�|�G���P��>/*n[��
��m/ �s�a+j�.�"�N��ǡ���Ӫ�[3S��cj�B����1F\�tsEVrH�]���1>ԍ�^Ou]]@�����[��åpOP4))�o����pT��i���~����`SSӨ6+��y���ݵ��|{s�r��( k'"	<�Dm�O@��БU�Mΐ���u} �ein~�'�T¦�J]�4��t�~��h�� �V��3�ǻx0X,�G����"��H�.�q�CF�y,��Àx[�?�c��>r233��Y������J$��0�X�]�(�Y�S2�0 t#0���V�%���E�4n�E�2����T���G�#5�Ͼ��?��'��TdT]���`���1�QD������
�Z�X��]M�2H���J�T�킮z~LD
��M����5��-e���^;d�mr�ɿ�.��JzU�B���ԼCJ���˿��p���]-P%�@+��]�9G���-C��%?)�(�"�nH�LY�g/~��wO��Y0�Ov{��{�/Ϲp��WC�ys:���:�mU��`���#G����7:PW�����?r����Ȋ�Ө��M�Ccݥ�[�5��| ��))(��u�Ƙ����-�eX��f�{��$ҩ'�2��1��J�srj�����zj�%�U��r��=��޺���YM��D_!�K��;�N�<<��Zn]}}��50���HaRS[Pԩ�q_��h�egow�ؒe�ae5"I��I������)��f�Aitv2L)g��ډ����}�o��"��u��1���$!�y�$�G��H���b�5S�]Y�M�íM�۷Gx{�nB[
�n�C�j���P�-��~�Cļ� 	���Mh#���[������ܹ��z	��Һ��M>��eVf2	[<@�Wij<522��5��R�y��{�@�цJ����z�F�E�8��@���?�,=�0��7�d�/MmN��cjA/;����2�hqG��S���J��>z��/����[ ze�� y(6�5��C8ڇ|0��s+T���S�k��������"c��ivP�@�g�.���N�s�n��;Mr+n�w���Nv`��z�'�٭w�r|�?����E�1_���Obr�7[1����#�۷o���& B�!
bu'�Y�<�DCMm�]� �6�st,��4��7���Ä�L�V��x\hZ@���˗S[�=.Wmpշ7N�tS���8����ٝT����6m�PV�M����ַ>�t�hɞ��j@�P�U?z��ᄀ���pj 4lq�{i$��CN8#d��X���Kʴ����Y;bKS���Cj�m��)����H�K&��>��[@+P�KO���H>Kk�@�s����!���o]��X����i�jԱZ�xxأ�.�B�CNK���DM���}�o��N�&�����13^��P4���d��}呚k��Aew�2���T�]�X���Dj	��+s�i�Fv�ͷ0�(����ଔz���������(�7+U=wK��(��?["��J��W�/Í��:B����w")�AF;�5�����J�,^��>�Vݠ�&��:��&'�ڮ��ȓh�T�K7e��k����Ԇ�<�ڣb]Yg����e��n#Mŗ��ًuwN>����^5�#+��.�8�x/GK5�uڢ�iӜ8'�v���m��2��ʴ�Mk)H�4���S9�&����w0 V@��,o�T������,|����$���:6��P3557����K=���yAs�[��qԽ(����kji�����zpȱ���J��.��~1h'��E���`wW&鸰z�ƓVVFb2ci����"����������kz&��s�[ȵ7�~��e�w����^ʳ�>/��� �� �B���&�TTa1N2�	���
66�������ή*i��Lbaaq���N�mjBX��~����Qp�YJ�}G��~�������xR����k���ׯ�y���"�yY�H';�L���2��L[988��z���/t�r�L#_�~���޲A���7�)�, �(�a��H��Xse췽�x �W�`�+��)�{{E���e�F}ikiYhyj�vȲ���7�t���j�&IpΔ]N �w�b�b\FZ�2)�_H�A��L��&�Z1��W	�-7>^P6x�FIz�G۫�/��VK|ЬGq$C��ec�z��v���
ɍ��Z rm�rRh�v�nm�M�h�˯�P�.�}(� PX���aڳNz����t�ŕ��2�
���?��2�Ҙ��^��2����j�;_t]c�Vbr�"�s��{��8:N�*��]E�[r�n!�9����"55n��ń��Yy�@陛��̚��g���,�����9�O�Bu.�C�Ά��I�$�I���z��6������n��D`HKD�.�� ����.�֩
���Ns�� ��V)�}{d
����tK�'[�k�x�+�4S[������*PN��w"�p�s�K1o�ۿ@����=�����Z�m6�����Y֝�7���E��L��ױuD���*h��>��અE� ��
4
����$�������h�g��Z�d$��u�'T���
l�Ҧ �ՑWs^n��cU�67��Ng�d!�L�5Ԑ(����<{="T̀D	wv�Ia�z�h⣃�1�p�*z��1G)�?al���8�F%�Ѵ��8���f�00�=�}�-""K=��+���k�xE>�G|���6�~��N�lh3�X�G�=mL�+B�l~��}��evv(�n�j�t����T,,,,���%�n���t�	1���7��X3g,�x94�Li�L� ہ���p��`6��L\F^�n�r�(	$�,p�jkh@M��ǘV6 ��\.L+;����4>��&�)�&�+Z���UUc�JO����6���l�� ��Dv�j�~��a`J׹�����?����~/�2��'j�M����Z��$5s��O��lc�4�!P�t�J���S���L@���h��a.�lZ��&��L�Z�88iXT�ӷ�E�S�p3��27�]����H�i(Jh���tV֝'����bL��:\:�L���w,�S���TTTȬ�"X)Q,{��0�
+�E�Z<���I��2�`J���o�t-�����P2?��i�U���"�0n�-)�![����� \��Ą]���M�6b�I�)4�n!U"��143;����XB��J�ejj��]`WK6�k_sች��WR��na2��#�#���0�5S��\�)��.S���a@ R9c��a�Q��`vww7L���\V��\���Yꠦ6���p�i?�ǎ7ͯ.���l�fں���J	�9�)|[Hi�����,�"��p ���e�(��?}���������2�00��I^��ؔ�W����WU��9!~օ�%Ւ���X"b �sT�����n�qw� �C
�k�ܜ�Dg�q0�d
���fT�Օi��u��)�*4���*p����� 3P\U��S$���6�J��a����S.�U���f��R� �.�����<g���^0��i���]��S�Z"��`)�B��d۠���D�*wF�#k����	� ih�2�7��MP�(=��F�a9�����TkI�7a^����f�Q��T �$��=��ʿ���m�����D���o ��q̏IèP��a�PM������=>�R��x���E���J�ؒX��\�2�M@�]pWq��2����Lʋ�O � HQ,��`i&=7�y˖-��f)�5.]r�K#�J�0v��r������W�hn�LII�#���55b&���->�����U#�0k~��+�Q$�uV���ٚX�+:��N��>gep#@y%$k�ǏgT�f�/@���9�@{́p�A�r��#j��j������x%%b[22������� ��%uu�Z�<�/d��c��DfZ�պ��-˿I/�j_:���JE��l���f*��t�����V��CϹ���=I�� �9ҌT���
h%���q�Tzf����3��5�o��7>��K�1�)82%(yN|���̀�ի��4J��]rJ�VCY�ꔔ�Ҭ�Ps���V�� �0zw>��=7�"��<e5�3u<Gr�a,������^~bDtG ;�?�829��R"�:��8fP�=Sc5������v@�]���K7��;����6�r��t����-\��0V�3@q�Z8<B��hqhhh��wS��m�N6<�[��Yz_�梁�_í�rҳU���%��ˬq�0�M~���Ĥ�S�=i��T0�N�ѻ�;������<�he� �����>1왮�eٜ��}�%*��o��%�aEg���x��T�P1��K����.dg��ڑ����.'��k�v�bM�o�Om1|�1��s���������R�3<����c�n�6d��I����Fl��JQPT,���|�3��s>���0�g�&o�4�h��秙p����d���X�����V0_Z�*����،��H�hA�D���΂���w��۾Yv9�˷�)2�8|�M8���.$�`g��Y�Lby����Υ&�����f�Xd��͎��ߟ���hLlF{�%T��a��1�_j��1u�c�ToqL���m�K��K6GY%Y?/��B�:-�;�y�^W��x��WeZeڢ�vxG�9�"�e0",��nT��5y��(��2LEؗ���QC��w%����1��O[,���Fs�M�S��j	���������F��[�����a��|����͛2-ڊ����؃^�$�.V��j��c��`A^̲C�㽕����������#��)������"@p���p�g��C{�2\O;}$�sN��d�d)#0���Z�?���RX��O'k=�ˇ�@RL���UKK�o]*�*�&��֥\*g�b��\�G؜����CK�T�C��:BRR,�}�'��u�j��'6��a��r�z��q�>ʂ����z��m���>���R�܋�|?�%QM�j�g�Z^�(+��㐿De�dZӗ/�����򳨑c2<����G#=.-�,��.�����@�e���VҲ43�?Y	C��"����mN��ab`�	��]��L���|I����Pؒ�����5]i&�Iꁵ9~��k���{|��^]C�Ǝ��J���>+�������)zyI�� -S�tN��L%n�����֝G�J��_љ�"��-����M�J�V�]֞��@�3�
f��I=9�?;��T��]d�1��(x�ºާ����U�N����R	Koa��3�L���Ց�����h�\����[i��ӳ��N���[̓���h�oh>���իW����M)��3���.d����R�"
�J��VV�ᄱ���|�������S��O>�:U�P�ѡ������#T_�����(��$��ob�� �Oc������p0(v�*�C>z ��S�-߄t-6�i�`f"Mp��&�,LU{E0B�#"��L���i�Z\S�g�3tr^QQ��"�!z]}pP����H��{��>�)0=kK씗�?�onn��͉�>�R߯�"��$,rW��)�.��R12�Yx[��o�fW�,�3�\R;L���4~�qgtt�ѣG��-�'|�2�������~___^A���ü��dӵА���E
���%��eZ��ӂ�ެ{������u���Ij;�C��s$F���5�7�,��$
n*bA�8W5��&'���rr�O�k�	j�DD�UOx��
&�UR@~Dx�T��JOW�����L�LYy�,���.��oE�����B�y����1	�a�J��/"�W�� c�{=���렄t�"ڎ�oǤ�i)~���0&�@�}������Rd�g3�Hi�Y����%��=?;{W��� UU����H����4������O�Y��e��{���U
�����VT"�&���&��h�����ՃW�ĸ�,�8���i@b+hWVY�?���:��Cg���������߿�cgy������5̣;gB�͹}�O�-4�i��7545�ה �ÏS5?;�Q����^7�5,���SO(*.>	Ѽm�L
�~c���f��B����k����>�lM'^P "ǥ�ӥk����D�s�	������8B@awτT�$;O"j�!nU�����*~E�4N�9� #6IUZY�j*jXu���Q4�f�b�ڈ�6�����Ϟ M#!!�Mz�4n�)b.#��LP2-�*�����5NI���rH8�2�wg��{ݐ���O�k"��s��J�N$�Tu��O���,p�9��GO�\�ؘ�职o�����s�;�kk^�sDn�dg7�v�O3O+�^\\��4rS+~�X��*.6���R.OWI��)�I���悮�/?ջU�?�,���֦TS�=C<o��뙹��W�?~�8U�*�N~#'�̮�IC]]�ʕ����g��]��J��5����Kt�F4O��@<�r����3�����1fM���>ȧV�,��SV;�ip;3�rB�>��%������Ԧ =(8X{�f��'��p�L�}��u���P:�f�QU���i3��S�)S	�7b�^F$���9iA�b�y�0�(����-�v��������m�?��������0�H���
��lS�MO7�ѣ4S�]� ��r��K��&A�x�t�޿iӦ #M`ZI�b�}����8<]��C��룁*�?-�!�Ѵ;��Ғ���/�¯߰ӥT��
�$ǝH��6f|R�}��eF��x@9$����L��c�v~�0 	�kKS9'���ܓ����{�!�8��һVݡPVQqP�6��! �U� ү����=�x�J���:6�8���
ŷw���aR�����ԚA���Ƕ$Eq��]��yKK���EEE�������������xq��	����MԲBBNk��v��D*R̈��W��ޙ����<�P^9�>���uu�ж�VR��+��	Dp�l r�[��)㌐h�_{�����\=�C���_����d%�C��!�:+G<��>�ߞj%�}{�s(;;;���ӓ����z�����ԡ&io+�'Y�������H������玄�C1#�� ��sr�ʍ�Q�#EћY8��ޗ��9T�ځk)�s�&D����8RU���U^VVXX(�9NP�O�1�755A�t��^���gv��wK�LrQ�Ӳ�����Х�6!{&�znn!l�����~H-?&��N�<����1I<�V~Ю=~��5J��s^k��F����j��vNR�����{�,'��e�ڇ���m_ߕ��@ٔ��ą_[%��|�u���ʍ ?���e��)�k��`e͕t��>] 1)��e``XW_�50x���$���<z�����±�k�C�}���f�oKBY�kX  .�ٶY<;�5�H��-!�^]=�`����x>��t�����/n&6��RV]]��ك?2F�o3�G�6�>#�VNNg�6^��&��#5p��&�~v� �>���?i�ʽw.��	�慄����:I��������@*�6�f흙�T�üm$��V��BR"{����6�&�B������4�b�萎�]$뱄sp8�뺟c�����y��<�s_���]��}������/Z�}�`$�8Ӌ�b�n8HZ���x��jV�ZB�B�$f����&Nv¡/2V��I&jn�p`P��l�V��c�(i��}�:tI�u�xAa�j�%ըY@�'V|~���a~X�d�ɿ�)��5���r��Iv�>��e˖(�m����c��}'0��n�A��yN��������ψ-��o�o�u�=��ْm�����8��>���5id�ΤC�{����K�'R�����h��X�V�3ˆƶ�S��~,a;*����{(�u�U���4�����Py8ef���nVz������==����?�8 _0���9i5��S���'&&>�3���nrWi��_���K�6��M�v9u[�nK���8�:;�0�g,�R��R��յ}��b�rM���;�-�לhѺ���z�ef���J6��Xl���fy�'�666G����#T��� ��&�������g���|6{�h�~M��;����R�w��B�4Z�@  >w�,��#	Uź�I�vj�5�y�z5<<��q����:S3�0��f���^P+�=�� �t'������AU���J�1�&��r,��*i��vv���iT��@�2��g�����vc&��w��3�T6���Ny2T>66Fw�R+�������EQ�-��ߎ�`WФ��!�K]]����Gj'�+{�˃؊����X۷oI��"��&VV��c�,��،����{f��Lm�]����R��S%�m�:456^����X�h]N��o5-*)n�25ՆB�D��v�\ڑ\o�O�D��ge�}���-��0'ҿ��N�B��M2�����;��} ���Wow ʄ.�e�am��k�8.Jm��l����u3�OQ8C�T�3=xv_���������ʌ<�@�/c��nx���(�]|r�����f�F��Ò�[6�0�̨��X�[h(z
>�V<+��p���3�l+%�y����g���ؑ��ST#v
���~۝1�ma-�A �9,({55�5i��.���5��?���a��
;��8ɚm߄?�(~����f��m]+����ג�&Fo��0ε/�{�uH��YyV��?��Ηa���7���Y��2��mtrr"
ǹ��iA�ܻ=~�s�Y+_��Q��㣘����['�p�@�]�wFY�&�9G� Q��ۉlH��n�dԍ(8��j�ؾ@Ȭ ��9U-]�^���h&)������S��ףYYX�OMM���8~7��l�~���Y��U�tOu�����L�x��!�k�[�M�B=9��l|�r�����_�R��Ԥm��7==�ʣ��Ԃ����;v�Αݾ}s���..۩���{��&�t��L��.ᄐ-�7d���Ǐ���\�&���[�BCCw�ݻw\|F��+���+��'F���>}��f�� dK���ZZ�����M�&���X��6�l�KJV��O�(�o���!�ܟ��S����-òb��{7�I������u>������|W�-��f��Op[y�����.,L��3�S����u�ЗPmQ�"<q��x�ν��[k�C{(R:v��t��ȹ�ؖJFE�������<pkE��������'����:��.BqyQo�'�X��x s�j>��u���ѝ�<����z���[C9����iCi����ᾀ�y��~~����ଐ*d������57�bM}��[�̋����'��NsF1���(*� )!)�5�U�P�Oo�el���@䫔�%Q�Gi�쁴E��B�>��ӊ����,���\��v������*))����Ԡg��!/���w�ާ[�^�r��ο?L��)P;!c�u��) %M�7Bо��]�_�|h>��S�y��<t��ϟ#-����[y��l���qډ�W��9V��bNYg��2̱0:�c��u��Q�s"���Xh
Lr�[��JF{�7E(�ǅ�.C��8;�6�A\] S;�� �v�]ٹV��7�v�3�^2V�h�� \�NZ u"6n;[[���:$kYq�(K
� W��*u���9� y�v�k�L��-j���y`���L�Ie���l�,VgM��F�=R�l�W�����i�Y���I���D��꾜�	�R��Tt��)3�� &8�f�'���h%( ?<�"���w$~hl<�v��9�U��?]<g{!��}H7���x�n7y������p��Ǐg@�T�{fA��.�^���)(q@��m�v)(�T��dL�u��1���Pzt���f�.*����=�K���] �&+����]k����޳g9���C��|{敶��	d�V�z�x�\e�=i��i�	�8�@7���Жܻ�&A|��Z?}
u�8�F����'��p>yAW�u7>>���$�[������~:8�����F��?����:X|@.��V�� ���>��j=,䊎} ��ay2릎�+��&�����Al�@�C�^i>~�x W�wU�r11������ؕ@~������P�ՇaD��0�p˅��ë��mV�UVB��o�lĉ�C�Tfϟ��8�mq������d�ȏy� ?<R�Y���F½{!�FG��������O5��SQq�*@p._0��88<�]nL��g�^��m<g蔯ع�}<��C�%�}�z�H�cU�O����v��HM�9O���q"�Dݱy̶���5��k��$({N��P�r�����\����ળ�����)+(W�#"#����4T"y͍N
M���(��W�]iS��k�o��������SM�1\�7�*���7O��O��a��Z��%�/���w�����.x�e��u�{��'졲 ����!��MUH2�J�ee{�{"B����wO�}BDB����䷝�=�q2��K@u�� -u��$)��3@< �s��?���)(��N*lĖ0��UhM�oR��'��IY����<���-C��޾�3���]"�����jh0"1��S�$�������+��u�[�����A��H�%I� ��/���Ќ�d��e)���/��+�Ml����#��(���B̢��5\�Z;s1nu �����������_kcc#4��(�2J(��
lQB��sM��B������Wp��I�]�A3�����is��'�k��C��4�|R�.��)���/_>���d��)�</��|A^�2�����*�+Q�vΥ-�\w~�'�[=p�g�sg�p�1ߞ�XұDMN�X1������ˤ|��P�����w�o�?���͒�[�
���j��]�D������B�=��7��[殺���P���?��o�K�|'!A&M�0�����>�9 ���s�)5�칧����W
�4h��A�zgGGi###���Y^�V���'Z~�A�R�w�=�ԥбu�� '�)ħ��Un���a~�֭d_��|S��^�9���C���Xjoo�fL}�_-!���.��O�*��]b��f`` �}0���+CjU���ҿ�f��nhI�{�r���K=��8YvN.���u��b����P����k�Q�TpU?��[�{���e�r����\�<�;��qTpg�	5xx��/�d	�����w �&&&px���y�C��$1`l�&\�ȉϮ�����nSH?RkKK��opŻ�]x�jk-�v����'�-�U��"�Jq����ɵ��~��]�eoȼ�-<9�c����P$pK�����PڡE��4gh�~c[ܵb��h��K�n>��������Ez�ڵ��g����[Ma)WU�4� �K]�Xߌ���C:Z�Aq���s	�o0�@���06���?}ؤT3L��o���+ZZne��v�
���FO7��Y��~��N%ԃ���y�j����q.�{�66t�>�^���mm;H��P�i���w� �]\W2��c�D�?���Ķ��E��C�ԃ�_�p-��ݽ��ҡʣ�Rf ʾB`xx��3e��frҷ"���gggg���y�����x&�խ������A���7}��Y���T�Ì95P�F��UQ�1ϗ��G��X�jUگ���������6����8��#��AT�?]S.+(+[\DJ���s�<�f��9x�ch2��O�/�gA��_f��qؤ�o]Od�AQ8�.̀"�*�i�I���*��
���LIU�SΝ`[�*@�Wc����ar&K�@P�1�>|8�����6��3�Fr
�ъ��}I���N�;�������㎊�5�s��Z~@e۳���K>�ؕ �Ѯ*�1?(O�)�b�B���r�Q�[{yɃa�����\-j-{}�F89wi�24���\.��;a{��`:�(�G�5Y���u��d�DF3ù�Om���ۄ�5�ɉ���:���@>��wt�'W�}�
�]`�˗/wd����]h[;�{aeݔ��\�g ]	�7����OL�(�/1�b�����4n��0UW�~b�����m�i��jrR	F�r��b���H|��a��ڙ`_ʇ��@��� D�YKHJ�*��5��슄Qw��[��d)�n���_/U��&�Ru%�K.�@���p&�5p���*�w9�@xd(�h�4�)��� $�#�}�W�.Ⱥ������mi��-IձM�m��Ȼ�$]]w e��X�PA̐"E�%#����v:'dfr�.��Ɩ� ��J�ob�� �Ҹ�q����(���LN�mk����_@���N�x�	�v�O��������>�J\Y򡇂9-���{�؀�Y>����#�����JY���t�8��Ą��}�p��m`bZOI�0Q��������=$���Y����۴�j{�^�.W�*\��AU�����4��ax����1|r�Ņ;�������MV�ώ� ������<;��d��� �E'����ӧ��=9�����.y[笠��
���Nô�{W�o��t2�	6����ND�S:ݒ� ��:���t�һ~����瞞�&3ї������^d@K(���F0� �<�m�j(���<�L�[���n�5#�1"�mK��u��^�����;r̝�֎Bp_@����秱 ����%""�K��3_�-�ժ� �}L�Н��[�:���3��UubG���~ZXx�t����
Z��nL�Jd#��!|q�To�z�8<鉌�f���R���>�(kTn\��m�1~n�;����e���wC�K
��
���\	�`v2\;mt���ӚA�V�O���������DuL����.U�{O��!��%$b���"���ܳ�ϟ?qL���p�V>?�@�_m(�̱ml#c�O�6�Ӏ����!�i(��;����Y,Ǚ�"!W1O9������3�ROs *��66���x�>d�,YEE�,|R���X���,q?DzI%����'>�Uu�$��s�������쟮j��d���P�!�Gvיִ�	,h� �@%AmR��6w`K%q*g�����k����4�3d����EOk� 2d� ��Y~Z��,�Ť.���bZ#!	��ӈy�l�J����4V�'�1��O��z�}��o$�J��#�����h1�,c+��)X�3����R�&a :Ys�/�pe�Ț�?��0��y{��-�����砦�Z�$A���4�c�ɡ3�xC#�]0�!_������ �4�2�i�e��N���U���9���j!� ��F!����!��>����Q2��|3L]���'@jڒ�� Oo�V>:35��_b��EAi�D���)�P���x+�W�Z�z<�v+=�چ�=�nBC����3�J"ԧ���3_�+;�H��wvn�w�m4�L�
f��� ��?���ѡ����ں=[���)l����^�v�H��4��,����95hB�9j{��" �TXI+[@�W��~�6�@��`�i�喰��ɦ"�	�wA�l�$R���ԟM�IU�*e��vZERJ�}g�z���w�b����9�o��ï�#���$p �d �
{��!M,��8Z�.p��=�����8(Z�E�~��{D戄L<kS���{�c��r���pi�]?�ɬ*nV����~$�}! S���TO��fPh˼ǝ�	��f�]O���i.}Z��0aU�Bs����k{��hU����;! L�<ht~UWg@]HEx!��8�b��FB�qR���i"�ʄ^]λ���CXBңlM��*&�!	s}	���Ɍ5b�_���	��xԊA�B�Ī���h'���*���;�,,�O��Y��f'�r�3N�g�^��O��/����ȭt� ��z��V��m��BWo������7��s�]�"�Un��_4���ׯk������̔���$����߆#���hM�Ђl�S�{��a)�Pѻ�~W����7{3k�hO�4��M~��A7��jTand�E��" �	:�l������p�G�h�㸋|�ր�߭���뙙��r���pÛ�ܓ����u�m���B0�dښ��t�0�\�����d��q��ʵ���x�S	�%}�\����e8��Fk�=UC>�,���U_�O#o��������b�ƍH]M䘷��	�fL���n:r��
q|�8_��P���*��Ʉ�$>�Y���Vr�[;r����(ܰm(-���¯<L��ʎ���E�]#Nd�y���6&��e��ŀ�?AM�f�/_��Q�)�]]���$N��A|�E""�޳���OG��ʷ�OzJ��fn�rhȵ9l0�X�f7t�1{{ϱi�}�]Ǩ+eePN9^�wj �d`q�b=y2�q5���3��a2Q,��ب�q,\���c!�o)�s���օm3ιw��v����,�����v8I�!���#��]���/��Z�<(�p�������)Q"2QxzH��8a$P�5W�E�&(����Js��k�&�ʹ��^��	��޽K�K�@:Q�@�eEǜqsۉ�=Zۧ�O�8�>�f��B�
!W�;��~���������t���L�K!j��kntm-;�xţ��K�^������!��ρ���eU��lz��B�nI߹�#F�.�#���ߗZF���E>�m�N� ro����ݛ�(:Na�fg2�w��f��;2��yʨ�9Z%"99����%M-��8���J����8��oX�pa�caS�=e�C�v �Z1�pP�T�&H��π���ϨMi��W���s@��c+�R"@�@�r	PPRZ�Z	{�8�/�]tf&����EWg���l'�ߤ�X�r6���NkL��O��oo�%���� ķ��s��S���^��i�v����|�����8�5�=���T'�����Uu�)::����l�X�
��]��e����嗀y���AZ��h��a���<��`Hdeq��=ggO(Օ�p�͙3�*[	*�jjk�!q�%[�V���Lyɇ|�Ɏw&7۬[����)@AEe�|tFom���{V�Z������>�����MćJNǝ�Q8�r���}�$j��n�z9�����m�Ǭ��+3+v}��_�3׸�U��j�s,j�"�"�C���0!��v������*+�X�`)ǋP� �4��7t6��Ђr��e�T��o���X�	�4a��=	p}�Z�57�:�R��H��8|�$T��SSSw)*;^� �����j�g��8"�M~�SRR:��k�R�$5<��#��5s�w|�����ޥ)�3�\	�g7�b����d�>/*@Sg�#Sm��S�i��8]8�70��Z�N쎗�=	�����8��x8F��"U+�,n����� Q��[	4���G�p�ٍ������M{���#u2�)ː�r�#v�����!ǎ��<���B�s����4�X�JY�%9��
v�l3۪�E�_ ���Z��	�uT���kϱ(_	�pO��,�c�.�*��4ྜ��$����P�,�� �Q��p�̅[ 9�`�����+� �]{��x#��	.����U:�F\<Y \��X��=��$����`���;⻁)"OT:����S��H!qj-���|Z����^�V�����遗��Rě��Y��o����9�g��\���EQ��k��$%�*kB��j�,�fL0�d,�a쁘�knl���lNtqv~�](BVR:E�8�yy~���{ÿ�����FqߟA)[�ؙx�F6�ő'KYJ������[�4�ݻ4���ň!��Q��P�׀Q_�h(u���k��9����n�sju%���������߹s5C?��T���w9;�b�2vO�币\5�"����'�{�4�q�_T���j��Ʌ����<xW���@�27�!ܰ�2���fj�՗/_�z�~=6G��wt����!����1��7{��#
T�i���c
e��t����"��HE+�MT]��BZYӼ�{{�].���Bu���N���$Q|��Wu��*�NUf�"�x��U�ȍ��{Q�7f�+�������5'�1�ٞt��"���A�)z��>�!ssz`� .u��%XOP�Y���z���rV�������߉F�}'��}[��Wc����#Qy���7��s۰xѢ����[yEv^{���E���I+�znn?��wab����WZf�:�*qK�G\�F��5�}��wAC;��-Z��3<����R��kr�6X5&��\K�l��G��GFܨr�@E�.=#���.}p�.55q$Q��@�y*H_��ĕ��]��d��nMMMA����g�����"l;;�N�5�i%9Drv�,�zP����Pb�A��2�1�J�(GjF����.�S���	�6�p���u�7��N���T���4�j�b���FQ��o/^īh�͘�"��[E�@��m�k�Y��~����X�h��W
��8������Qltܒ�3��>���-Q���t��h�F�ZPY֔�n��	[�b�D����ڎ���Hq�~�.
DP���֐�ҥp�ƞ='�o���!<�o�eq���̕H���q����{��B:N���c�&��mj�	�Ŵ��I��]��}��]�Ꚑv%3Qh�9j�D��t�O\8�%IEsS%28}���k)�p�~M�T2�r�G�Jx���,�یՉ*ӑ}oWj�Ml�!rr���zAb����x�x�;4�C�A8�9RQ�7Q�Bn2o�L}���9c���ca��O49����mC]2ؘ�M���m'��t�C:���G!�\N3T�իSSS%>Ö��&1�	j�I��\��gPt���*��F $�GU�=��Vq:_��Ã��:��m��x��t�Gƪy����_����q�im7��Ӻ�J�o�k��|{f���d���ݻ}�
H�4��(�#�}|�� hi��0/�U%i@���������])� �����f����>�]$&��*���j�7
���AK�B�K}=����gFP.�"�;��f�T����f��WVV٣�E�7��k�.���6Ȝ�é��K�8E_���s��J�䁒�s/"�N~�K]?hݦcK����p��9?�%?�߿62B�D��?}�
���y��P�AD�⡇�-��n'�ɓQ.h	�]��
�m�J���6im�o�ݚW��^���㟗ѳ_�0#������A��s�o���̞��>�5t�w�ܑ�@�12u'.�ӡ����p"�d����DBY>l_:���-̷�#n�y�;Ed��l�sJ���|�v^* p�RP��(S��9�c�ri�#�4����5��x^�£JԒ`O��VT�t����l�F��V�G@è����j�i	��������$YP :O���]��bRL���7lW�e�Z#fstH��*n�CzJ��u�&��3��7�𗊦"Ui���)H ��|{ �zV`�8�*��4��xw�
��gLŋK:��߼�����-X�ҿ4Q�..6�&��г�����vws��:��mIT�[v$j:KԦk�>C/��3�#�T����QAȡ0���X����'�_UU)���f5��3�%�3{����H��"�fRd���f�;	�����������}@�귔ym�{߸zu�ڵ�!zZ�����/�s�՝Ri8��uɒ%��xqhf���-�6�VM]V�z��MGp��f������Ȕ����|*�����g����+：�	�P2L�3+ܙ����dfŪ�/�T�`���\鬔��?!PxfZԦ��?"����K
��qp��q"5�!,�L5U�����66:(�ɉ�Z1"���9�EDp�a���~+"c/oy��hNy�1�6���;i�ˁHhN�����O�d�,ߔ[0��<��� �ɿ�>����A����l�BQ��������Dko�����CBu<&;إ�aɓk�v@[٥�n�}���)����c�%]�J#��Z�ۚ8�hZ�����O
�è�~;;L��`���B�C�pjQ�;jMq#>))r����2!LM���.�<��]8N[���5�F
E��!e���*|�.UU|*z�2}��<�{��J�'{Ī9����79��B�Ju�k��chGmB�l��Z����(����]k�l CaE��)>.�?+Û�-!�o�Z!ur�5y�3CЫ�5��H������
E$�n����g�k��Ar7	R�U���h7�'�R33������h":����rMJ�=���9ei��R���p(�z5H�U	z�Mėr [�KC�F��n��(�}��ɓ�.��u���Y�TB�!��	���~`F�
:�f��i�WD���|> �օy^��K�.�X�i(Y.��$WQ�5��F oh���*2�tHi3O��65��/��%����{�?~�Hɉk�:�>�q�m�H���1U���z�\�u���� v�&�M�FI��X��u� g���5h���5��q�9~���Sb}�����B}CH��[�d��/�q��&U+�@�p��gIj�)\���:��)V��*�ѱER�"N�E�5~���d�_���{�Se�����K]����=�uߑ��'�v�-9�ä�N�c�Z�۷�����-�� ��}�sM��H�󑓱�a�D	IL��Lq;���PBth�+�S��s'>>�U;n�u��t��3�����h{��MЎ_:���Dʽ9�V�-X'V˨a-���+��k4h���c�Q��	�.�<��s��q"6�D��S��."Nq�%El�MG��c���K�����Bh��Y�q�UҥF�8x�ࢨ�`��]��6	��<߈駨ج�A$�Pх� �w>�3'�?�%]�BBǸ�݋�����/G�����(����v3�5@]���D��G��G2a4�56����
��񧥥|��q���з�
-k�c�MNN�/ŀ�Ƈ�@~h�n'�����.�X�Z���]2,��z�Ğ����\��#Q(�dddn�>�&8#u^�ג���?�J�����1�T]_���w��s�O���� �7oR6�b�����^'�:��N�Z��#�P���LЭ�ˬ���.�.M�n�o�d����b��EkW��n�����a7oB�����.,#Mu�08���8Fpd�C,k~όq"���5@�T�Q���Ή���knlhh�>}�����$�(h溺��ˣ��6\�2��4u�l���6��h�o��%wsA��&�N�f�s	��PK���V'2�̈ ����.�G�)v+ձ�\%�r�&p�8����Sff'�����ֻ��5���3����p�����C��J�{�q���֖�sr�!��	�T"K��(qN!Hve�i���0V�����ܾ����G'�����)a�o�Z����G������&�T⿨�����~�������U`	��U.�8j=a׮�x-c^L��Ν?��ݻ��혣�xn����b5v�����X������wD����'ף-H+�o�Ɨ!�3(x$�Y�.����6���f�����R���R�;����CC����Ū�S牐��{�������sr^e�Ƞ�|f5փ�j��������fq�[��R��ǖ�gMґ�ܾ��?4�StŷX�Cm\�g�|������	�|���Th���}vz""_��&9����aj�)R���b<��>C?�x_n�j�s�b�24 l�0 �T�L�Ω�w�T@�'�G^�+O���-���^����kD��{#�����>�G�@�-�t��X88����~��5B�q��_�6���kB���>|� ���@VW��I�^ F)�j��HJh$�y�U�JR\:��a����B����5N_l���J5R3Հ
�O������?�����2Nx?r�������(ť��t߀�N,}'��p�xg��VXJ��=���Q��~�dv���lE�QE�TG\�]�@�&E<�E�֯_o�J�[;Z-�xj�9�RZ�7ć������G�l1�z�nS��7�j,^��H��a�z=|�.�tH�:��D\��e�޺uKU�e����M���#Y�����+�.�gB͘�iv�Ӝ[�&gM�3`<��[[[I	y�K��k,��3�_���'�j�u���Z[-?��:�M��|݋���+4u��j?"d��S��	m�.Lp#�u	�˸��}jj*τ%��]T���˺u��恎C��k�*��^N���S��N�ݱ�\�i6WxѲ�GDQHR�	n�|�D@;�`:��|�c!X��V8wy��O~� �]�o�ћ�i��U�����[C!�͔P�n�kǋW�4!B�bi�x��̤���=����nʭ���6+>A���&1/��9��EB0��;pI�{�r��}A�P�e$�Ɂs�f8}%<����O���i��+�/Bb-d�v��W91��9�����!P��
�F�k��l<������"!	]-.>�ok������'?��j/#I�>xff�xF�[�.�DC:��S���t(.��Ҳ���+Ҭ+��{�#��0q�bݿ�wW�LU2�u�ĉс\��y«���E� .�t�F�X�&�fdfZ��L~�]��KA�Ҙ ��klFi��0���&��b�`�ڜ;����>0��f���!||�CO�:��@�[V������o�i�43df$�<�E%2;;'���㩄Tp��W̦#3�<���qF]H�6Z�{V�1���!s�s ��#Q���R�_�L��e�\����(� �(20�8)(+qr�p2�����QF��ܻ^�/��2�4�vp�J�4T�� ��}y�X8I��0
��������E��Һ:::.!�V5m���'����Em��j�ά���B"�ԺS�j@QUf�	�s[e Y!$d�Pږ|�߆:�
�3�<�1�5��BVy��u囲k��� �#fꚔ�p�*d��V�D�к���cۻ$�9��M��sP����q��#��[ը�L��1(���m�S�J��&)�Vk��L:���Z�=�x��27��i���		ھ������H��\��ƾr�J�95 r������J3�>45]7�bq�xYV������ގ�ڕ*Y^`�|"C�%v�ŋ��aЌ/?�I��,���(�K�koV7�t�fq����K�'z1N^��_�K�T�)�?�(��}N0�ZLl��d|�#T"��ŋ#��4cl���D%&�swB.q�F텲p�
0����(OP���״��m�g��c�������j�T�[��w�_��N�$�
xZ^��u���V�Nb���!]}}���QA�,��9-h�F�%�`�Bf�$��  q�S��7{��<����e.�לhUz~s�Tw,�RU��JHU��}6��l&�_ ��ԩSWKKK�R�;�;'<3Z�����Sl�� ��vT �D4x�6?&��2޵sgm��V(��==�O���C�|��C#��g�eC����ތGH����9A��Uf� �c!p�-n,Y��W��2��V�������
 q�~3�z߽;�F�~	�L����q�rn�j�鬉�wB�kK�R���2������(�l��_T�*?��C.ke�5���$��ZZ ���p����1u������^uj�R��Z{��tv��L�)����M��<�'S�|�#4��7C0�dی����8Q�W�v,8�����ƍ�b��p�zzb�r)�io�Pl��
݊�c�C���I������>�R)h��!�� �����T���c4���DՁG/�}iE�S��Ӎ�\�_AV�f�L���qsۉ��l�����$̰�0�%��I��k�UEZ�!�+�2hm%@�}�;�[��oܹ Ҥw��cv�={6oh{���Z"2�^r���@	:::d)/5������C�A����
������
�(C�mp�yfz w׾}M�Uh]9���~�	d�q
c�~�^�M8cS�7fg�WA���&�(�����z'�B���ljr�s��ZZ�	D�ײ!����7���<<�d�`<�-�.�~#�t�#���p8��sA�`��k��<b�?�1Հ>���!	]EX����"U��a&�V-�T�pǕ�_inq5����ߓ����Ɋ�n�T�F�ڵ��n�Ƥ�\�q���n�,hQSU�cz��-m`"ll�*��}
�3�v@A�^��v/��>�d�d��G�E�{�����LN�%�����(��~qI�b�C"�N@(�/�d�������jM��)�z�.��ڬγ��%˾�jxy�F����C�7��ǥ�����V$>j��$O�Xy�rlOg�����Ws�s��J��{b�9������5Į�F��v�D��Dل�KL� h`|�3e�ЭsVH<'����Av�"	�j����;^��Ƶ�a�	|�	G~~��=�0ҟ?Y�,�.7����Xd;��MCN�K²�2�/��n�A����3�s_��J��J8��Ͼ�3��gB��u6�S�RL���ԙcW'ck��m���Y�d�k���� ���B��Y�f�R��99� 8�U˄6�n�$sy����X��7q���FZ�-��A�Q`�"܋�Rt��n�x������@��M��D�P�b���%K����� H�5A��ɪ��Y�|)ܞ♅yG-ɵ�l�'� �_���3*��3q�i~��nE�Z����%�xd	�[� O��-�Į�����U畗�u�����Z�Bk��r@w�7n��n�읗쑨;��5:�������f��6] �7˘�N������Υ �L%�M]B�v|�������BSUn�p&�ckk8�O�D�q�:��퉻�*ב��2�M����:>���
7���"����7�"�?CB
�mM�]\PL&%EA'\= ����FҡJ-���h�׌�:kW��mW�nI�X憸q9+�2�j�qI���,��d�gB�0QWiE��_��� �6�A�ٽ�hv.�2��j</oT��9�2���Ep�o�1�匰�	���О,���TE�#�LB)GN��������M$�BO셸�P�6�x�1mI�Ԟ8����)�ە��j�����)3��S�Rd�Q��p�3��Q��W8��iǯ�-����&U��8ea��-(��ړ�Í��׬�2Sr���5�+��y�H�L�܈N/]#��f���?�Rջ��L�)(���ڀ�q%�(�c����<ɤv#���t��|(��A)�R�$��T�F���ف�5�6�~c8�"�� �$��u�4��u
��'\�����N�7$�y�������E�)W&�py
�Q#�V"�U�4N䎿!I�Y�����E���d� |����xr^H4��w�5�Z2!����u��i8��<��ׅ�o��F�����'��\=r��%!�Q x��M�pG9�7�W��Ȱ̭�H�b�~���^P�-/�b�ƍ��s��x��wB�#ʶ
	���@�:�N���ϡ���ȴ�������m�ۄ�,k�X�?��F���N��<wF:aNkn"&5ۧ�m�Kh�Ϟ}����ˊ�Q��z[���h4Y�!1�Z�B�ş������o���,E��E)e���.Њp<�z�9�O�	��60�"鮉=p'�)�`@M��Z$��1�@�wB�q����߄=p���9I�<jg��X��z _[��s�O���x�h�dh����ʃ��!YYA-�r����9�+��X������
ߧU�4� 111��{A(1B���c�0B�3=�Us����A%�Rhx�b�L��.A_���R>����Xx8�SjN<q�`8�W�}��Bכ1<+�?���>�hH��՞�{�O��7m�������&&�W��(�oO�g�����f��c�<�U����fѫW��s�*F��<����1m���N���������C�U?~gQ�k�ѭ�孠�C�m�"�����*Jp�a��[��7�ڰ�g(J����M�%��V�kN�G~�����S�L�y'��lM�h���I�t������.b�}i���h�F��T���絽����G�|�hAǽ��/A_�8��ʖ-[D�^��2e}��Ny�ʰ���!��???f~�����t��~��2r ��1����Fg#�,�Xgu�V3WZ�pm�$\�w5e����i�A�F������o�4��f��	xe��)��A�L��(t�2O������{�1�%���eH)b�e��\����N�ŋ_�^p�kw=��K_��pN���Cp�eXX؁ȱ���z�V�L�̚ǜ�����H���57%�>;�����3zV���E����GF�����.���3�6�ˁ�����H�_�Z_X��(R+˘I��i|Q���a81��B����r�w����}<g�Q��e��{��}9��љ|�0H��U]"ɇ-��1��uk���)��d_�;��׽�C�>���⪏��37�jErU�I��]����67p?~<3�-f���ha�|%h-��gJ���V�J�,P���+
l+M_}����-�m:*�l��#�XAk��l�<T�zµyLdWz�r���
x$몒V��A�6�[�����gV������q'��-P���	�K�� �ٓJ��Y0�+m��L+�~M�������KbO|i����2vqi����'n;+]�ƳVY&������{��r��Kǥ�������[R1?e�G�}�����ܜE��?���d˂�P\j3�P3<�'/�4g[;/��Sz��x�!��'�`���3��C,�y|u��WNY�����ȭc����������6+�hȾ_�'?��?�P��3����2���ZN�W��
�D�@���}������V_I��3 �C��> �`aԙ�k׭;!����:���K�}�&��{������T���4E�E�	��*�[��ݺ'��m[ن;b}*%Z!۲��_���lZV7�U�⿵{���ѹ��K
���1/�#_qt�=��i�������S�K|�z$S�}{�O7g��6T��gܪ4��,-������_��}����eDF��v�G)B/Q%���֢�ۅ�!ML#� h�;VZ��ip텠 	f���5�c*wӏƍ,E�|�vZ�t��6������n��ILZ_�CZ}�}���e���E)�8 	�������^Tu�m��V���~VV@ℊ~��F���m|��@Gq���X� bҵ�d�����o���ɋE�i�\��d����^��)��߀j���2⒒�` j�*VU�{��x��e=�G7�z�sQc���;զ�A�e_T�S�$J@�>��ߴi�s�7L�)�Y!���_����z�x�JNWWO��ae�c�(����Q͹Q��d���a�1h����|hy2:x'�-�K'g��%�uRz�s�>��+�����c���)�6�šϑU���KB����CT�]�ee��â�AU��Bշ�tO �AL��y�ZU���
�8�v#*�X"5�/�	��lVCC�9�ut������'>�{��9`�cR��ѽ�oa���B����V���ϣj������ ��Bc�Q�H���,�9�Ue>�%�Ӝ=��q5� �t�X�0�C8��7�����Omz�ۜ�2��5�d7/�a��/���XYl�#P%2c����b����P:O&�!��b�Sqf��T	r|�Q}CCC�ݥ���-I/ܰt20Y����m��(���H1곹�������GfŮ}\N�XqMk��xBR%eee=S���6{��g�c֩[�	��lᘊ����#�������cd�����%�5{����5�͚��Y�l��
��Ȫ	�
x.S�Ͷ掎���9WW=$�9���B�h��<��!���!N������H�U��-������h���ր�D(eF��?�\2?�%��Ӟ�����j-�AZD]�r�4�>'����b�'�d�f�ɓ���X��_�8)��XWTT�ɯm�������z�}j�М���:���¥߄����t��珏��c�x,�/�1�9V|�m5 �)O��*4սr�"�5W�
�
9�������WN��wԷ«/��58������[ /х���׿���*9E�pߩ�]��c�����O��ޘ���~B����De~����S ����9������YOy�L##O�HJ���H��g��Y�,qnn k`Ph���..$�I��XƌF��U�0�<�G�8A�E&�z.�c��1����p��c�9{tO�ٳ���N�}�
r�{�����r�fP����~i�ˢ������~|�67�"Lc��7o�$���]�]o!�6"xϝ�0nsP`{A����P���W�1A���GG�~`gg7��0�Я"ө�����5;'��M���+{9;�#��VO�ܧѧ4��?p�n~��%ɸ�  �]݉;���l�>��\�U;̏)Ļ�s�⺔�jk��g�s�|VE@�����غT-� ��wo����c|����+�q:m��� ����Qq�!��X|͛U��R�8���rx.��5�J��~}do��y�"�c#h�{{=4���P� k7��\��4�����g���$�X�ӷ����q)"�m��C�Q�v��#9t�{ 8$$��IA���ƛ]�ܔC5Qy��JX���o�ud��h*t2��X� ��鯥ش��'	�%�ss��xA 5�����-���ܛ9z�;������c".~~��EdF$u'�_�#w�Ki�{�o@���'����kM�~���t���é)� >����V�f�1	�/��I��ҩ��g^�U�y?6�O���u�I�)�O?��
�?ܽ�f�E�Ϋ���
K���C��G���L--!I"�,z~��)T�L���:�;^{�Z03��6T����[��d�}�����p���i)�3�f���䕕��3�%���@7�u�V�"U*
��/�?:��i�ZJ�������0��t�2;`��i*TMb{u��/�ʔ�5�?�U���Te9@�UE��ҁ^^^�jN1�
T�mmm�H�P�-���0���{Z˼t~��'�r��c`�N�81=T>\PQQ�3�Y�֭wP�Ba{����a�,d�caS�~��7�T��g�]}�\ܾ�_�a��`c� 
����e�Sy


��C�8+�1ؕ��9A�\=4�f��n�Y��bv匜W��%c1���H3X�Rs��㍣�`��j��}��V����;���w��2����V���V:lN�%Q��RQ���19��Oٲ�!$!4&�!��(E���`0���<����P����������_�l�������������� ��tu	��M�j9=9=33���F��?է(2*9�C�F� �A	C���[5.��Θ��vd��?_f�}���f
����*�U^ً|w��}�w��'e���*��4����weҎVz�8xTI�y�zd�9Pe�AUƹOh�R^z�I?�3�-���4�� _�ŗb�?��xb�
q*jƠ�41���UWGq�ψ՚z�'00�TJ!̆��1c�Ur�A�J$7k�7�«�C��xj��U�'��Q�6��-�toA(�����Ը^%��I)�Y_OO2Հw5g2�Vr�'�*�ׯ�C����j���m�74ըI��.�3�T�Ȍt�X�I4�[n�H��_}h���h���
vZΝ2�������+���m>~~t�&�úk���uq{9`�Y{��C�������A<�mm�=а $�F���Ǐi.��!Q���������<
��.�<!���aRS�������L��R`�a�8nա�lY!��(�m����-Q���Q�U��BX
�Z��%�@���RZE��R�՛Y�_��Ga2�ȥ��rroBNp��w��,(���y�	�B��Z�D��>�?��I
�(���u[*H��}�US��]�������*�GJ,��N�<8�Z�z��2�����fK��|3����Ej�FY҇�G�G	��	d`���R�b��y�!�[�1�x�NUj�Z��y�'���9q�2�UP ��H�*4x|��άf���8@|�Ai�Q�l�i]�؂�f)��ԃf]I�xz>�;y}��Ǒ-kx�����6N��Of2��f�kv��d�k�A��r Q��Z�������B��zȂ�Ѓ�7�6���
�"�Zi.�e������Ku��K�.�c�X�h[K`���ONNV�d� � G�f�Չ^�<���`���p��� ��䙠��s�/���e���H� R�h����%$�0�N�����b@a�W� 8t��v��s��(�����@U�L�����8 �U��C_ݙzR-�x!�2J+Xʳ�!�'ԽE�|#,�)��Z ����~!>)!�2iot-ѧ"�e'۬)m����0Z0['2� ��]���j7k�KQ���j���ՏQ��,��;'TBJ�E5\H�`K:nd�_J�U	��}�Ŷ$PL����(�(j��%4�'�v ���(��s�k���P��?&A :C%���>}Zߖ\j����\y�2�Zmmm3�Y�FY�N�C2�TaSס�C� n>%�5����*p]of��������n�V�:��ф�ڪ�Z�¡� �<xpx�>��/�P�-����wC't�h�Bm��J,�R+q�$�
��Lp�({��-a��enn��&2����G��گD�_���ylU����t ��@��sh�������<�������bb�5Q��J��}uq����s��N�}����3�"Б�ѧ�:Zeh¥��6!�}�H韯e ��P ��<��R~˪��i_�F<�ؤ�~��i������2jc��TZ�-�������P��~��L����a��O�8 5�S�F�ŝvS%UU�`֠ܬ: f��N�R���d�]�B�����N̨�h��׍��6�Y5��x'Zw�X� {����e��o�n ��}��]�!X�s1쭲��/c�/�+(E�:��o���u:�6��t���4��&��3
E�x�)$���D强��k?[YE� ���@kL͍�&���4ܵ�݅����D,�WPȆ.A�B��c����F��F:�Ç���H�,��L@4�9�zS���C>�Gj����[���.��{���7o�xg��m:	J����jU��X��P:��{�O����s�?�EB�@���k��}fFZ���*
����A� ~b?Y�ȇr�M���Z�AYu����Yn۶Q� �,4̤6��9C����W�`��U-����{�S��+���r<�D�rz~0a1P�CY3f�م�H뻄k����9����)�����˒|�6�d6=7�=�vXkσ��gV��sj"���^�j�{~;+��5h�V(����D�lNe���J<��1C�%��ܩ�����2��RQ�]�Zv��ս��SuŌ��v[+ެ��L�ooGLS])�l�̞m�s�nDD��'y/<��f�/L�^�����?3ܐ��|��ͤ�w����D.)�w�����X5��nr`��ީ��p�n���ǪJ�KÑ��Y�DL�`���_-9��795���۷7cpW����6�?VI�g��H:**j?��V�%��Ol�y]����h�����"u###�ih�|d���2�����	�1cjH��U�^�sYs]9
�T�C�{��ڵS '���~�V� pn�c8D��k��J��ܳ�"� �nܸ87~P���:0��6��Y���2T64P�l�����`՘���m"�ܞ��&�ƧK�!Ս����/�srJ�	@�;����U����5P:1"���tM��g!�Ŧaˌ���/���el�/ P\��zzH�iq�����1T�ݭ���GF>�XE�������j���PN���V�0���y�NE�2޽�|���if^~�������Ix6#��`������.�a�7����tF�x¿��q���:�%>��t�1@�D#]S�R��b�jhp=��Y�q�RՇ@� ����8��<T8�|@`4X��k\^yy����3�P'����g������r�-����fb��J��:���g�G���0O�@��͛��.��bOOd<����Xg=����'�w��:8)\y��пM�B�;4:M$�ڴ���vp�$;c���]]}��x'��|��!J�#ǃ>!t��҂�����=8-�d�B����+ ]ez��>�u���.\�h"S����!�C��9�P!I��m閖��r�s��~Y�u��<�֣f�����	�Pq�|ɜ��/n��V�U�=�yt����b������}4c��C��.�.������ԡ�L��(�2߿+�vCVJ
\���v���Gw��mW�jy`g���Ή��GP��i�[�kxT�U�h3�H!�L��9��J��3��?'���8wz>�z�޽7�2�9��n\)�<�n��S��!sݱs�_�?�_� ��!w``���q�.��T�7��D��[*ξ�	�mu7�>�)�%�{w���H���`�+._L�� ��C�|!g[�'��N2��'y��ݿ����ͭ��>���؃tAX���Ha�0����M)ĉ�����%�}���-m8
aL$"r+IO���-[�0'�::�J�zWP�Z�5k�ق�����Y:rO9�F�@
uDH#j�3�P#bX`ú��=H���ڴ�D��Y���-�Zr���d��/����X�����S�������YK��!��1NHHׅ@+�D��T`���d^)��ƣ�/u���j��ﳜ�y�YU/��B�O���s�r��ٳgU��y[��>�=,sh	vuׅ����2.!�4aAc��r�� U�*���=1Y��'9� a?�{E�y'v��3[[JKKwg}P�Z�'=��s,�i��UK������s.)$�zY~�u�8a�X�n���H~�5e$��f3b��T�j�� 7L�����V�m�<��אg~uź�@YF8�|_��L�����@:������{��kG��f�Y��b�b0%je	k�^��Eꭍ9������P��QŴ�������ڋ�����g����Y�莬�2�(�-ح666���d68AlwMX嘛.1��� ���!�ckk����%�����8?�X���`L��!A��1�~��A���ȷkG�	 /�X.A,j0vR}=�X�,�O�n�۫&)�n�:���ܻ���\]���D"����|�]�8k@��T�����ذJoϠ�*9_R�~�E�;_?�!!�md��	֬}I� �@`�J��/���S�'q�V:��>��R7�b����.NN�7n�P �����܌��IzO胕7���V�!�{%6ԕ��W�=�� mR��pSj��/@�!�_�<
Z� �t�f�*|�0$�R� ��\ɦ��RZFF�����v��ȡt����5 �e����<�H�V$}*����c�b}�,m4mp�z��D�M/��UB���3Y�?���� �������{��*;Ҝ���4�;-llH]X?Li��7a������w3.����I���T3��q��u��*���g"aMI�ǻ�&ءz�,v���?Ӟ�h�����iƹs��f2�K�8��`�� �I�X/�y�r<��З��'i�A���i�^���{Xfa�I<-˸)UՏ��r� n�,��$�Dי�f�`9>V1&E�����%���مN�ȸ���$��/d��������226Ʒ�=����d��쬳��)$d��{_�; ���Xh�D���Ҏ�4�`�-OD��w��b�R�=�h�>�p���'����� 3&&���p�;[~)ZS�ӱ����.q�ϫ�Ӆ�42օ�b�۞����/B��YSs��e����]�<=�8��q��C�����w�ۭ_c��o֯�9>B�>���U����ps����G��.$�xA�ө�oL���U�^lJ�,�`���ަ'�΂ȓ��3��mDl(G*���q�J����R���Q��ʠ4�q��*���h2��^�`s���wW���*�Xl|�}�Aμ���d�����J�fy���3Y%y���Wa�??���a�s�H<T��*�`���މ=�K����K�3H�������q��j{>�+�#��d��С*��J8�:�"J{�[N�Ò94�9; I1����&��BAqh�W��JKWN8�b���eX�ѵ�S�x:� g���;��q����Ȇ���v�ٱu�&�+a��q�Y�T��J�kԁ�BƷoO��}�Ť�R��fł ��C~Ph;��	-F�����7or���t|SG�b�/����"m�5dk��)Dݩ���k�9T�'���cqk�#��*!ZJ��e3t�|@��E��[�=�(��4�T�CMرc��݃�� 2�|�7���E-���T~�/|��R�P��lg��3E�)&:z�3��E�lW����?�IZU>U��AC�?+k_!l�j�����R�'�.�Z>|��#����0�G������dƹ�Ϲ׻g{Br�O�y����
���:P�f��o�'�������]�'��b��\���"�Zݽ�9G��=TS[���C���:[�I,���ܼ	��W���!6k0]�!W�27x�ÁͿ�ִ���N9Ě�ۊ�({'|�ECaH�:�����,$ࣨ�Ekkk	�\�0m������	4�Vk��^_gW�D�(����c�̅q]!�O�z<�x�?���~-;��@@_��2�B0X�5���z����o�9�^\��� d��8������ �E+i���mRx�B�Ň���=7���/��>QlHc|HX���6�l�[&=�L�>C�v�gZ-�P?JnѤ~������dr�UB����n���� G���k+��xv�}T�,,,|�ZWW�����]�ڑ��N��ǟ�8;��s�κՔ����q"o�h�䓳�}������
e: E�BP��i�Xա	�r��~�@퍕����n��<'��#�W�@JJ
}���.��l�Z��H�h��E��v����	v�*믑U?Y�lŪ��㥥��9�
�*n��#B!�EP�wf��ː8�2&�!*A.N��^�1�	z8�K/�Ď�b)(F��b�� ��M�=m��F�yK�j�����-�k� ��N���x\����-;4�C,���[�d��=ˮ���pK�U�5�f��ҕ�̀�G,���.;����'dO^�{b��e�1��Re��!s�6����G��I4����<��LW�����V�=��� B���Xd}�|�Ԑ���;�����{��5����W��߃Q��KKK5	��*��פ�]�l��o>���X\[iW���܄-�������^����s<D1j3�0M�鱏#~���'~��2��^<�d�1�-n��G;B(faaa�A�*�	nS{3��,s/�A�khh���xx�b�W��1�@d�X�E?wt$�Q����1��GV����,���'�������k�m����o~�F��H�\�G����>��O��6��8�ߑ�H�3�}�nD��{�~N��[D�~5/W�Sx�5r)XChg�b�����g(ꉎ�oO��sW,�5��6/0�ӥ�X�0h�ֿУ{�3Bػ�W�2�Gw��[��P�ʟ@�=��V�ZݱL��5k �
 y/!��	�g{u�A�����'Z���ީ=Q�^X����"S33���["���wN ���Zk���E���"�������t@�Wϋ�J݈ׅn�2^�}Z,��W���t�9ͲJ��D��%���������ݻw�U�	�����tuu������
~�~����G�s�����ld_�ku��L}���o���>�g�E����633�6)��\�o�M��E�ʗVZ&l��s�I%���N":�0��"fR{f�O��La�Y_���z��D6o޼�Mz��&�N�����CO8��+����9�����Q��-q9r�)|��ʭ�g?dCqA6o�mnLa�%\V��g�r�^r)xնg�'����$H>����L�ӷ�E�#N �������EF�;����}� >����v��}���w�=��F�D��ps����(����udĘ��]*��x��Z�/�5H�aA�3r�QJ���V��X��{�h8~*�U�jY5c��=.�����<>����T�|G����U���jڋ*(pvs��X�h�����L`���!!V��Qn�QM���g�El�z ��En"���*?�1�{��4��z��D�w'�l�/#��)��R\�C����
�;!�m��yV��I��s�~&j� cdu�@��C��֫j��[<�W�'�>9�rҷ��(�7o��<���<w��	$��2 ����"������J{rrU��_��oA�d�<�r�I��F[[[^N�:T��i'["��"kb������n�Yw���P�`�[�+��&�?�{
/�����j�w��As�wt�+j~%ux�5���y��V����kv=�~w�pb	���4�g�E�똕�R�Ђ�,�~�wYt9���W��DI�TM�TU��p�p�����!<��~�H}��e�w<
�Cd1`)� �,<l��{�� � �x����BV]��0Pom��0!5Ig���ɚ����E�M$��h#S-�]0�o�z�J�h0�z��CD�C)�J�p�U�������PD�P��HF��6ke��@�̺mdg�o��h��fTYc��Ǣj�[/X��1�hWr��U�&�<�z��Z�KHHH���`$O�?�~�u7ci)��/�?V+��}(�cZ�]
hP���OC]�z�ָ1Pmt�a��Har	�6�gѦm�喋���8�ѽ�N�^��o�2���Ntf��h!��
� �/J�P�����Hm��m����j�W^��+�j �j�v�)S1#�y����U�'�ܷ��}[�) ���}�����l��i��DQ�ט���i��]�M��ˊ3�]S�5�Dc��������Onn����9�' �PO�R�V�w�� �o+E]����8�����ё6q�� x ��@|`o�W��i���n�x��<�P�>d�+��HK���̜��3�ޥ�Z������Y�!6�8(�����M�p���(��Nf'?��טzR�FGP��c�<'����S�&���Θ�4Ͱ����n���C6�Ц�QSx:��D��n�'�f��g7�K�K�$G~�N{���jdf���������^���������(m���Z�?�VTO��yE�	D��&�����l�/��%r��-~fU����O ���@Zm��w�&�T2��^8#DH�M0�[*���6��{E^AŃ���sm�:n�U^���������b����t~���C�(�3��?�M����+���%!.^��� �(��_<���O����|8'd1��:��5hb�W/Cֺ��u� ����9�R��;vm�SDj��C=�:T�n�(���A�4:a�Q�<�C���K���zj�"�l���)��y�M�/$�iCK��E�0�D�yB�����(ӷ�!����^8�EKK�(���24�>s߀��dv� �et�ֈ���ef�M:�.8��Hµ�,bN�����ߣɱdK	��P�YYA��u��g\e��JJs|�Q��#i���#�3�t�j���M������!�!����м��Z�M�i��ƹ��Ad[I�ʃ�� ̅�\ɡ��T�w>��h��R4T��ԙs]��X�4�M/+f;!��1�	�\���Ѓ��v,����E���\�֝u���Z���~[��~�*�<r�:��	����Ӆ�����6�-��p�v��`�?{�)�����߾m��%�z�u�w�����O�oX+1ao���H����ȍ��ڪ.�z�7��&c͆*>݌%��痑�/�z������h臦������Mb�!�惛'^�4�D�GT�P����+gS����A�o�$��փ~��l��4_�nUY}t4��H�UM�ު�Ws����&#��G1!��K]읱�(��x�u�f�y3�Kc��v�4����􁹹��uW�v��3����g4����sX����?8�0��~�H��L&�Ҙ�g��)�qZ� (��1�N
����=��,I���(����tx#���ӳ�	Ǿu�*YD �C���-��IYC/�MOK;P���ӿ'�TFN�f������y£��s�W����K��eOx�B��ҟU�Vꌗ����#}&p���]#RSS+g;\hR���	��&�t�cb�/�(>��ǝ:C�z ����Ü���̕{d59>�F_l�����4��B=�y��������|||^���x�E���Β��_�&��s�_/�J=�k�ܮM�1aj�r�7���'v��"�+k]S�����o�3��ծ��JTsI�~ɚ��%��r �0=��5g���^����� e�
I���R�I�'c^��s�)[B����՛�zì��MSJ������W:��9g��aUUՀ��"j������sZ��Tا��0�O���Ŧfff
	[]JiD��Ѹ�՗Q9ŢBB���4a$�Gi����Gw��]���	D�a���O79[��dg\wm�u�8��vO���̇�A��v����W/=p�m�������h~������Yb�X�5��p|����w���N��G9a�}5S��� i��e7<=��}�v�K�|NN��1�ʪ�D��`��3��۵��q8\d-ȣ@\wv&��\9�<���� {�v�L�[��Y���&&vj"�2��������0&&�	Qi�P��tгN�#8+�r��t��gyy�]��c8�|$�ʠ˝�*�ڞ�ե�$�<�� �G���$?tuu�����*���Nyy �!�yyg�H�g6?�ņYk.W`�)�°#{Y�/U��,���7�B�j�7ʊ��SS�R����#�]]��k˗ao9!>��=��DVu�}��2�<���3�&ǿV�Y٠L��f&�u�b��+2�y2|TR����dݭ��:�����~i�K5���RVR�'� �{��-Qa�Y���Y�	��Z<�;�{��0��g�q�~�����,�Aat�`���չ*`%	�9�L�+
��U ���D�T�#P��X��/t�6��V�&.9�\�����Pl>0`_l���j,�L�f�"uФ �ج5:�$�{4��8<�ٸ]�Ѯ%�n՟�p����Z�}"s�=r��������9�Ο��^x�����t�������H�~s��@�ol�(p>�6  G���Ȱ���Y<�D/��d2�<6}�����[��(�oe�`�9ͺ9�uZ8ժRC6?� YȆ�+N~�2�2���l~��i~��|��W���\&���@Y�ϓf�lbe���2�>��6Cs/��,TV����Q�.�ΙO�'Qx
��s����/�;��x�5ZV��fk1 6�E�d0�`"1��Pk�0�� ���)����X��3:xi!�����NO�@�������A��e)�U�N������+�����[ ���JP9?�+I��	G=Yݏd�kznU����������?vK��nx"ܰЏ�K�޿#R䐷��9��^��7_SI��K�V~���Ð��pU7��`]�İ���|Pĝ0�x�N�����&&�q����Se��3�HE�A:���,>5�W'�x��?��i�h_�Pd�������<�Jq;h���~폘�GA�PVV���Q�LN恐��籶9�F�b}�7�>��R����[}e���m{}݆1�*���*GQ\!�q�Hw�HYjwh�5��H�)�[�a�ҵ��u�>;�����\�&���:�#�˃Yo���z�L�>5���s�9�B
��t"�����ow�l�1B&�#ȡ�.w������@g�)+Rn��`��n�K���a"��:TK�S1�)j��x�)�:�Ͼ���c4��I�kUz唬���T�0�!��,.�*SH�-J�6�'���@�候@��ݒ2���WI�761��OL�i�,X��5�⡒?��Y��0��1�ẹ�����H�300�
L~}��9 �t&��h�/�mw-�A�E42s�&�j�$�M�{��J�|ͺ�"Qa\�)�\��"�i~�W�Gps�|��EP������ērR�>l8�x��������)��KƱa�uC
��h��&&H\�"�����ף7����f'�@�_7d������s�R�bBNr�a���-�O���]L������Ǐ�5�3�0u�w�P�n1�>�Z� �@��Q�[�$�ngJ�|K��Yʆ��P1K�x=VV|�۠��<k�֌�Ӊ��8R��  r��v�����hbz�Fg�4�3��[<k#I���[ϵL�:1"��Xу�I��Z:���ųeIN� !h��kgn��6�oO��+#+RR�=��������`��<�X�ؕ�����	��u���E]��>f�@Y�m����9�މ��yA�.|�z��[�}��.����>g'�L�g�bD�xS6q��-M􉕕��2O���ńLM�+�xA�����W �;���8��<+�Y�ҟ�T���a=�e,��~�"��P���?n:v�H:L���f��N͠�Q~y��$����G��I��Ned�, ��1��Yk@0#A�i��/���ksvr���Ҍ��F�����h��be��^]�0�:�3r��B>Vj"����V��1<`���fW~�]��T�� ��I+#���㮞�j��C����#�SGRX���b,�#�	`$�� ��r�f�e���Nj���	��MJ�{�/����㶗�<��ڂ�ܷ�ʹZJ���%~(Z����H`���$$$���#�mM�ϐ��Rԏ�\�5�����]��߲�&S'&�F�q.�����|���q�!�5�ަ��2=��#c7����qT� ;�{?).���n֝Ɛ�-�ܘG�<����w��2Z<�,����ط��H-�`Cl���5��1��3���e�Ȏ7��q�����!ͅ���v�'��l>:hLٗ�Y�OL�}�G�xғG�0Ca��1fC�B0nҐ�sԟw�7T���.�&�����x�GpۦG�w����t(��a�Y����*];u�W1�K8�+s�44�ꯇn��i=;�
+�ۯ��l�Lm`���IX<�����`j�5	����ԉ\C������&��D�z�S�Me;�%�AC��:y�*z���dc�$jT�E��yJ|���y�85�tTg-cb�.��T�&?~\�����M���)�u���b�L`j�kB^^�%��I���9T����ҳ�e�o�=Y��'�����5i���a����9aERVW�oo7_`��qݨA����(�]�>;c��k#�n19U�p�0�;����KVrv��J���~�h�Z�j�9���N�g�a�}�����Bl2��N4�Ѷ�?n�u�����8���z�#s"߰.z5�e�j�:�.��l��~��ݚ��	\��J�a����̀�Wt��S��{�|����zN�c$8\� _-|j���GO�ʙ���;L�����.P+����L=mP�;�&Qg��^+����?W`[�����M(..��AU�?��|�fG�-P��.0`��o�r~��� d��e6�>x�w^䪻�bIl�Q��|�%�e���C�(	�M72ʌa�ȁr���P�$Wy.�[�k�2E�����ى�B�|To�j���˞Rw��_��+�b�����6&-�95\��d�,�	�~{�0�;F?�I	�\^�{C��Fs�i~��G���[^�\!��摵-�1|��l��C�Ŗ%���&L��u�~�$��Ur�S�Y��-{޶�sݨ�����hV2�R
�����؃>���ц�-k����6N�����{��kHeW����&�n��
��JX6C���V��D��j���uW$�����L`YZo�'Ž�d��y�w�r����4O�JBI58��WtQZ�;�/[>f��ivb���?�h[�8�Xk���R1�pv{'�VTA�nl�4�׽�J-W� ��cc�]c({�䁫E� ��������1��Qd6B�l,�ຓ���Fjj*�{�m�:�-��uU .-�B���^>�q��
��R�o'C��B��Aڡ����3]zG$4t�õ��Cd#r���qsϡ1�k��컫כ(o�re_8�E���_�c��A�*+)�F��(L�ԫ���0�o�Qv)�i �����k�Efmnn�|�t��A���fX��n-$w�:��'��P,�e�i��������v+�LI(��{�� s��w�-�A��	!����#�]T׾YU*�Ys�� Z�?}Ux$?�������[Lo\�W�L��z�ԅ�.*��?�HD�� �~gU��e����j__�6_r� �Sq���,W����8<Z	���D�b^@�����d��T�s<���K�N�%���B�Z�W���8u�hJ}�K#I��V�\N�G�B&ygl҂SM�1�"�Q;^���l�����T�Y���0�Vn��G�-ϩ(�4BJ�
�s�կ
?�[7����Rq�Yߝk���R?~V@����1�0��v+�:�u\B��Ϝ�u�ѨP��PS&!����>����^݆�������K9���u�!MV#Θ��C\o�4��@F�!�Ԛ�L_��Dy�����=��j;��ֱ�u�4)��!�,^��� �Ӣ�:��f��� K�7��~��@�� �.�.W�=i���狭ь�AY�cv�p��&~.ed٭\�z�<|)@�H &�D��yj딇F��\��dbA�l��w$�l�z�^�b���Z��iA�e6/��N�������iC��oΎ��-F)v?O'��o1�V�SI���Ԉ�&܋�#
��j��	�:�浺��f��`�b��ߘ���V.��Z �����P��L���5�d1�$٠7���*�&'����!ӄ��.���I�Sf>Q$��V���cE�?���8���B��un�U_OOO��dc��<!$_Q�;�Hz�"67���3�0�>>>0dE})�&�Fс�*z�Z,��}[��D���э�"����a0Ôt��(�\{�Bb|��~i����X,��{�K�0�>,6(~�aܢ���:����b�;������-�r�vf�PQ��[?����g��H1�	�Y������!�3�����y;2�C�.�r�K��h����&	�K8�ŀ��Kȕ��K�`F�Q��6ZH���&��-��ie-�K���e#�1^�7
.x��ƈ.�[~������f���^��Toe�3�>Y�j��At`k<,�qB���t�٥��^��r��p����櫪��>��|ɤ����;�WZ�.������:�̍���d���NO����zK�Sb�{=��1D�2��K˱��n�/�h4L�R�z�3�9�0?�B[6�]�/r�����@�̵��9��!��;ɲ3O�},�U?��&�Ɗ�����f����B���e<=�4�������z��=��3�4�����`G��T��Q��N�ݣ4������]<Z��<��@H�[ɚ%��N։5�`��w[ͤp_�ȁ�Y�N���p�B�%�)��	��/�d�[�:Ƨ�+2=�� ���%��Γ&��8D�|%Q�y��H@3��#K˨��m^�$a�j����۷�e���j� �87a�?)!f$�* u������xc�����Z*�1�Sv�_�';OsF�N,l���S�Aff&�-�>צH�"p���e���	1����cZ�8iG��X  ?���$ѥ;Gݗ�Ks���xU���h}�n���E���$�Ђ:�z�v��~�������W�H�3��>��/8���&#���qw� 8��-_�Y/Fa�7�Td\��n����l�`��ͣ��������l.��� ߘ��Y|r_���.�4�K
F=_��X'��W�3�Q� �n"�܃%!>tQ�E�l9N���F�)�/��4���M'������x�����w��x��3G�ƀ����v����y+Z ���b��k�b<�Lt��(?�5yƗˇ����/(z&s��y �ԔӨ�@�uC��F�\�����\��%Y�$I;��?5�[K<���Q��a)}����~E���}\{��=uMp���^|����-�h#u���6���q�K�Tu�{#�dJ=?a#M�4�\�&�9����O�0�܇�۹�c��Ų��R	��.ץ|�6���AP%*>OL����b�sK
��ƹJ��v��ɽ��!Gre<�vC^�����Tb��h������\|�J��H%y����j$6�Y�v���4���'j�[��` 3u��4===��F���[�+#��Ej"3�Q$U��2`$��EB�U3�ѿf[J_��m�)���eaˆ�/��fX�=�HM�0k,W�L,@6�)¿0a��Ś��9a,�z���cf�ឣ�^I�',;@-������"�A���k+
�k�`3N��IAUY
�[�\,��Q��/)V4(�ߴ�fi۞�[���
�j�Z�w��{�^��~�� ���¹��k:�`�n��9|���o�y���Ԩ�G��|��0����K��O�D�����1�P�C���H�+�T>�jE
��UM��i*�5�S�l�3\�����b����'c��!�v9�Z�A�!� ;���'������/��Ҋ�1u&]Ⱦ��Hx&�ekE��S�͞?.
ױ�	�S�� �r��~�c��C��8p��:~��P��vlk��W�����|Þ���{i���>{~f0��u�s?-��B���ϼ7���5h��@u�[`U�D��Ba2(�}�
�-�\��9SD�3CS��%�w6�t�,O�P5��s���J�{7���ŗd�}�<�� ��g��Z�Ref3�Ni���R����U�.��ʣu�8d�XzGuW w!��|��ʔ|�D4��s��!�p�N��]�;�w�k�0	�cMw�_������͈ل�O����;�����3)�qj��zH(�w�p:��ڱ���~%�r���Nmc�Rt�bL0��}�^#݃��[h�:s�'?�ԟ<��0��/>��Z�3��A)��
x ���{���y9�D.�;�X��E7߃�~��m�"Yu�q%���w�?��2]�7z��|ȏY����0�J��9���:T����s���	%���u�%&�f��I7�qO]5n�3;F'��4ߤ�w"<�k~�]kjh��}��c��G�R�p_�:E��}�����-��-\��O�x$��zc6t��#��wgR��H�Xk�F��}�0SFhEڬ�˞Ho��~�$<�L��+A�Jc�i~z�3�e�1l+��yz��Y�d"��rZ�2�1�D�z�^w�V�K����_�t� 9��1���v>�g��CC�@j��� �p3��Φ97g�:C�;�X�&��R1H	�Jk�zr���+��@����G����R������ y.eV���֟|���?��}�g/�j�m��]?���d0Fal�c��e�P#���2�vy�����v�lj�"�D8��BN$��0���l:��x�𽷊����ja�\X�|��~5��A�%��C��A�W�p��I1I��%��-�sy(J9�r ���HpB�b�K��M�[��'�ո���dwL-�ֲe�ز�];u_�*h�!�)��M~�֐tġ���+0j�U��kE��q��.��c��#�_��twu���ƸI�;��	�j*
�Θ3d�ko�Z�IZ�h!�n�H.,�Mj_o
�T�����5H��
��w{�-pq�5��o8z���_Q� �����>�x*�A�l��$��i*@ق�r�1Y�;1w0Q�j!2C!um��e���R���Y/�fd�
�Wm.�h�h���V�H��� �O��a�������TG���@X���WF\s�WL hN�G})H#��W1Z;���j|��R����)��k�JY@�7��K��pb�|;g t�9�L3�/W��g����i�Ɍk�-�9��;"Q��6��M���?3d?[0�b�0��
���`����&<O<N�ӁQ�%AĹYw���V���y6G��z'���v�hf�$Cf���l����_�����I(���g���HOҗ��3����� �����=חH�bm/i�>=yTW��p��J=��;�?8W��V��c�wq*���m��[;�Ԓ�!�)�FWA����C8���\oL�v�r��s��u*F|�=�e�8�ɮ��5�IԏQ�7#_^x��B�P�HL�#�틘fÅ6AG�<}����l� �+�����QYj3�����>�v^ߩ�ły1m8�F��Pl>;;{���	巻& ���	���X��
y~���I9�B#���bS*5��:$�p��H"���F��������ݱ���B�.͋{@}����亦�Pz#$�B��H��'ǔ�֎�?��V�.��=����]�x�(�ȴp�h��5��Y
�p1�7O�[DXxs%����9XÐ䓢ƒ�M��ߐ��3̓ѐ��Q��l�ch�}�e*�\C(
)n��a�1QL�n�d�+�`c:!��<��n�L��9��ׯ�ӻ�����	�~���&��#J�&�o/z���A"�"��ul�'cWLmJp 3],��*}D:޳�[Ik����]j����{�.��F&�=���Mf�v��vx'��)�SV���J���F�.�sM��f��0M�p2�l���p��D��]��e�:3��(ٙf���Da:7��;iQ����ِ��(��P��=K�`Z�,Q�����/���፵j���П���7�l�l�}1���ۑZ����g(��w�t����p�H��>v	

��%�£h4k�맹�N��#��#Ғ�� ��9f�X_	��`�Rwi�U�9����)mo)s51����D�&e��e��̗���U�Z\La����mq~�,n�Z�{��6�n�ǹ�[���ϙ߸�ȝ��� �n]˽����SnO���> �o�]���]���]���]���]���]���]�_�|�6������$*	=؁qA�ڽ�ՃE����S��}�(����}�鍸 �5>]O<��^9�X׷�r�Ӵ"���S�CgB�>.?\饪w��N��3T�͒OoM�%��A]/x!V����EmE������n���o�o[Ł����ԼZDD�,��� !,��c��!��%ߌЃnTgt�\l접�bB��*!ʾ�jj��?�;ܘm�����=�.FvL�O�>=7c$5����Cʣ��&������4Fy�0���q�����za�3��ɰv�Ԡ
uji�~�W�ƴ���ٞ@�y������kI٩z����T��6r��_��G��<�/�D�+�Z~����]�]�OClC�go���?}O�.��L�~6h[��ݒ4÷��Eb��ٱ�'?���E�/�ut���5����c��u?ߔGƞړ�޽{��UR���
]?U�PK`:&.Hs�~Xj��9B����@�����3�����x�Y\��]�������~��av�ҋ����&�7:z�h��߼<U΋���y���x��b�޵�\X����KW����3qu��UT򚚚���������(�bm
���n�õ��C����277��pUEⰒң��K����+�z�߃JZ-Je˖,��[R��e�E�˾d�-WFH��k��%	I�-�l1!ː��s����<���^w�|��,��}�9�s��Ae���P	q�"�Sm'�Dp׋0Aѷ�d0��V������o��AwL�C�S��?ݽ�\�2rKȤTĭE�:����A����OOO�\���b���H>��l�o߿��GO[������0�KPRR�-�ū^�RB�Zf�R���u=	�7�m"''w&if�/k�� ǈCǴ����zk>~������gҳI��A_�p�ب�Ěw��.G�����߭<+�u�����/�^�#���>�%����=������0e�9vqЏ2m�=c�NZ�5�r8@�����P�
�ء-�d0�\�GOO�R������~mӊ.���[ξ�fX[ض��J\������f-�D���� ���x�b��EN��G�^�4u�������$����<UO;�'<�70J���X{��s��vN����uҹ�
ї[H�~�ܑ詟��e�%�`�}u5��{O֩Li���*�[{K6�q��4U�W�C����*�����W��OSjB,M�[�����6*A������ס_9��)V�R�s*��ކuuu�5�5&B1Ȩ�%���Mۋ�0�4��)�K��9t��ԔQߌS	�#�f"�oF�������9���"�Z��_�1�7�S��ÿG�r3���{z�0pȦߦ�˯�x����՟��Ԥd��1ͦ\�>�[l��ۅ._IҼ~��QLLڭ[�b��s�;��<���Os�;K ���W���'?%��mZ9:�����Ν3%C��}łvN�02;Kij��!:W�4�ɹ!!!LE%�㏻	��=-�G����34�a�`7u9;�Y1�Y���-J���C�FvtD�hK�zt����e�r��a�
�9}����EuJ�9%����af�/���)��ߍ�������?_=���6^Pݘ���'�^���]����n�O\+د��s�<���+�y��G>������s�P���TEԇ��#�`\�ͮe���׻�SVj6� �Sl�̞]�|�Z #2��o_#<%"�Ã���p],��m*/��o�'�c�dÙ�
GG��ч2��^镕��϶xj�@��(����KН�8��3��TxC�NݺS�RP�{�M܄�<:Č������{�><:�d����!'���zq���L�˶~*��  ���"�ɰ "}�'Ff���|FFƜ�1Ew���ulm3.����֏������c-�̳�ۄ��^�PZ�?�x@�?�xb��]�\�KE�K�_D'��Ss(O�'U�_����2�?�IO���x=�������	U|a���#�vU��~;���o��;���f�����Ь 
Q��ݯ4�T�M�1��k��S�~�C���n�W91�)]䁮�Y�۷����`VT�O��1�r�-6 }�Q���R��,��2��1ְi+�}^U*�H��C�/^����g�G��t�;RK�%jh.�u��ۊE���*���C��o��ej�����",Gp�O=����7*�xT���xt�!�z����͹2i~�F�S&<f||�_Pp�����M^���%W�Ʌ]]�>�	��D_G,@�2�n��[���jd�E���q�/�6EP��X��:��^�3��Z2$H�UoP[�q���; "�����g�͍�2��� D��_�;���}�SQy��f8t�&��m:R��c*�f-E���u��|]Tx�KCA����!' �jk����MP������ڈ�u�o��l����|������U��Tk�+���8;
�H��\��^�s��1�YL��/��~�J�@DWb��׍���ff�k�1���]��y��mtf&77�	,#�������ʢ/!���)efh=g������u[������2��.�<���h����ľ�)���r���N@-t��w�P�X�|�����9�n�\Zm43'�v�jiY�c�(8E��� �y��`�ݡu��Vp��Z�����"�W�nQ#�cߕ�u�@��NY9Z=M�pc��vt�%X��dP�B8`����-Kkv����;<��ia���o��r��1��@Wt��s���[G|�N!߳9�ξ�<ۙ�"\'-�'T!� xu �m�v��$�hyʔ�0Q4詈��n3?5ڽ�����7n�*�gj���y��ׅ�Nx��hu���k�sKE
�.g�XB�Ɡn|s9�U�g`+���.����a�� ���ƅ	��Ww�m}���'15tW`^��}�X�}(kk7;;:ҫ�QR�K���n\;�:�F���������/�սx썅frrrܓ'�ַ�&Z�Ey�j���4W�S�������þ����/D��.�Qd ����|ɣa�-r��v��Ma�r���@̽�7Z-�7��yV毙㓼��|1�'�Sҗ�-3�=��x�����\C��߷��G_6�V`����l�9/�b�?���swͺ$
V�mK:��@(� !!�g���J"�����<�"����2Z����ILX[z���`#�`���j�>|��@4Ǽ���e��3�K+����	ɚ�>��FI����"�6/��oss�h�Wq8�xˢt���<�VN��@`�u�������f�#bbx`��>�P%�F�[�0�zu���ΐ��C��$%xfT̖�X[[㺶p���S�@\V��ֱNDWG'���>Uf*��m�\��!��[=�#.P����]��kij�x�cܹ�chȹ9cž;�S�fU�2n�~�/��˪.ʹWn�`Ƃ޼��jm��=�oz��DRaz
^&1V=��rp=2��[�<�v!�t8̼��1��n{r�}h]Ry�4����E[`��f�^��萙�L�9���^�:��][�nr���<���ﯧgf�
=�^@�u����4[��d]�Ƃ�Ү"�����M�^y�cv|r��Q8/?�?�sK~aa�2@���坌v���i�[��p�}�.��N�XM�j3c\�z\w��a�`:::�:���������tM��m�gb?�>��*��@�So��{�n5Ё/+e�+Qw�>��·���ʁ�������-���K�~���9�)N+�-{j�l���I���U����*&FF���[޲������4��@�-'�t��Y�fyKƕ�jE/(H&��֛�������f�h�8% �!����D����<o;��Fƌ�\�X�;1.N��U�,���(B��`�-���2��I��y�ec��ⱸ���#Q���!�&�(a��vaqQ4������z�G�~�omj G;�\6�D�+P"�rM�mM�v� ��޽υ�U�;���W�;��O�)�K��)|������5��X�#.� ��XD0���ã �`PX�?u�ĕ{W���rTהn4�㺶���#����^y�>�챩�F F���^��~��!N|�k���!�p+��tu�ZFF��tu55-T�D3�>6󔳅$�L�\������?����(kgi����~��~)9b�(��B�K�����\U��������\��Fط�0�����ۨq]Ŏ��D�聦-�w���<���'GA�gܥ;{z�SS���7O_�YZg���*d�ˇqW�i���*\wx�(R�>�M��4˫^'��!�����L�2oq����Ϲ�ПF�ݣ�H\GGw�����"XYi�n�u-�ބL-p�*�Ou�o�	�!,&��g{0v��j���3��!Q
�C,ӓ��X҃\��H;7D0I�&�˭b���)HcY���tP��+d�Rs�<g��w8#���R _J2J��Չx\�6��]ۖ8 m�l�j:@|���]\ǻ�S�JJw@L	�跈�A��H�8<�{�T�c���G)�-3}���Kc���͸.AQ� �wݨ���m��}v��A�rsZ�s�46^����J��|���f�++�@���Գ���PQ��~�����������E#}����AVJJ}A� 8;t�`) �E.����qܔ����?4X�d�;1q�B�٨0�b��lw��mW�|@!���o1�G-+3���h���"���,!I/^p��;�	O��51��v��zZ5�3o:�b�@,j���ڧ�&X߯�xН�*&ff{ �����Owi���K�Ʒ�mx��L�\��%�)',��������`�龜��3SSm^Ջ���,�N��:^����[��u��a�������%٩q V�J�X�>�ڗ���� ��@L�xdxi��`KT����}}}��^k<Z�ʝl`棄n�,��8:�N��Sc�?�u�	��o��n>������������6��ي9y�#��)w��r��B��~���&+Q虁�F8�_�(��wW.��RПEc�F�2j�bT�砏P�W��M���,�]�X�cg�k��r�G�=��錴B�'Z�/���Y��i�`v~���#�'��`FJ\���|vv��Jȩ�f��t~�6��G���DX:�΅�-�v~:�( �Z�ā��N�T����3%s��J�f��3�
(�2h^C�qFt#kl���-��̜N5������z���1�S��rZMU�:t�*C!�ʓ�z��ǂ�HWt5𾢒���n�2�Dg�i�R#O��>�EJ���Ci�K�m���e��։�P�ah�ro��r������u�f\����>7�SAy�����??`�� E��[�$m �i80�A�|�����;ڝ�?�����%�]cc�s�N%�}}H���Q��KӐ<�^Y�!�9UL�m�\=����QVP�dm�"���C�G�764��>���}ud:���̬,=-�羰B�C�P2�~�����D���\SRV����;�Ae!~���Z_t���:�����*��}Ŏ:��S��}�}�x���<�����{�����$i�<������8v��K��A�ij����Т������A�f���q4L�ʉ��\�_�.�32b	�����bj�]��8�4��w�V� z�����b+�sl[��@��9:�yxY{P� +�D�W�e��j��`��� B�u;:V���&����a<Y&��v�O��h~�-DA�Ģ()�����eTV�?���d�%�ŏg|'bm�.���3}%Y/��D� J�u����Z46��|(ӐH�R�ulA1(��н� ^�N�gA3mϾP�g���r~ˆ҇���5gff2��+�^�{���а9R�t�@��gt���9dl��w������'C(q��<3'g&D�Ԗ1�$���A��
dٲ�����}�ƺ�r�g�No�<9��w�m�$�Nw��K� 4���{�ߥ���J%//{223c���wSy��S�fa���'<�ݿ!����َ5�|ǁrbȭ`��oߞ��3��(q05��[��X޽gOYx7�X�)fţ�q_��\��}%���g@� l��{�I�+5�5C@L����f����o7��BPfTT`�Z�LDCd�����:��a�9!fd�����@��_�t��lȀ��&�T��ۂqK�;��#\�������;u�������-���I�%mmZ��e��N���v�����������V:�}�LU��ւ�Ru��7��Ԡ����3�a�*%` p��;&)@��?���RRlM�CVEE_{���q�4���MHA�k��y��F�����v*�V��n��k�m�m�٫i���'�JO�2Tݫ��?�=J���e���wͣ�,�E�z!c�yx6��//�j\+���]*]���DHx�XU;�Vw���W����g�\5��S����5���D��K�uE �T n�q�a�D|t7�*����R�o�e>�0��TP3H�B �{�-䒌 y������4�y%%2^�)*19X,6
���F����tHH����]Y:�z���y=��Mx� )����e��v�h�7Mtp=�M�w�V�gpJڇ�'�*5H�n���9�Y1�.$�/ !B��R�J���4�j$���{�>'��뺹�>)̦���������<��Fju"��/p8���..�����H��[���7�AYlq�6JW�	��������>�V�j���z���V�
�I��v������q��||m�3}@E�M9�����L���bd��A���Y`���e?�Yii=jjjBO��:�2}{�<��n�������[��-�	�BLM��@�`��Y�2`�qq��Ӏ{ cs�?�`�����5��h�2�l�[�.{�O9���AAA\ǖM�km���3[6ɑ ��-,,��-,,0������c�~=B�.~�\l�r7��+�ˁ�PJ�R�`�6=ݎ��q��4�ǆ�(���Ye��}��Gd%+�w�v�!���?�}U!=ݏ�!J�-�wn��+)��WS%d��^
�ۑ|��=oԭ�t:�Z\𲷲zWby�.�8یG���m����������t@���,���(�g�Tf(O�<���rGo�� �Xp���)�����/�A�֕�����Wa"�}K�����#.=�E�%���?f-��R�u���>d�_jS.�,��{VnU_Ymhn��j8ߣ��(�l Ef?^�m�KK��/]����˶������ܹ����%K��	ʱɫ�繒��� � �!��h�U4���a),tc���2�R�������u� fɱmx1��� �+��@c(��ڟ�]�G<�K�A�l����V���(Kxߑ;�hJ��T(�ر/���}{���#�hJ���!��!�W���,�3�����J���oƺm\o��#!�ϻ%��V*��FB9��(f�Z���֕g^�\1�D�� �|�v3��C�=	,c�tX-ԁ��SP�j�
<�s�G7�:::7.��3�lw�a
?��u���t�I~�ϋ�@ׯ�	�p)Cw�\�bŷ
�:���i4\����S�L�����7�m�I~)���P��$AQپ��mhh����Hc�����wL?Ozݸ�
�#�A�2T��de=����]��[����T<�ܴ�]��[�>d�AK��'��z"-#uW���"e
?{��? ����x�"�͡U(A�T����������6�C[XE8�X�R2�TQ����ܺM,6�Ύi9�h�10�s��.�n���׮�|i���+#Sfz����EH㕡@�T�TR\�{2���_ܴ���]����{�ǧ��x�������SSZ�	���A�����Ɵ�b�S��߽zS^E����{���v�O�$>�&e�HC��F�� ��a�~C�gh&I� ���8X��_y�S�)*h-#�Ɛ�,���B�)~�B����_��H�BҞ�6����E
��
���A�gfj���oqc�S3 b�6��(�25��H� D+�@�Mjk����_�Ʒ�c"PQ�<g���44���732*{>�/�(d^�}��rJ:�>J=����ֶ]�0؇OX�����P�y�����Z���t߀�\TH�cnn�DK<�!'��r���7�S�1L��q���ݒ�-�Z;Tm�����=�o�7��E"䙱13��0����J�� ��������IOI�^<Q\M�K*~�;{������oz�����K� �_=O��m�(&�ދ���D1.� ���7��hq����4��!��Qd"�l���o���`�Rs)3�-v�G���}�_H;c����������j��\f^^k{9~d����^>^=�cu��9�B���vԘ;p7�ʲ`�X �܏Z���-��<��;���߇��9�20`�q��^��=�G�[Z[K�����sXԋ��h����P{9��d�xbX�(rDjj��)M�J�B+��IvW/�\�����Ȟ���>`�M����_	�НW3�j�YRҽ��Ъ��Uo��,., ��_e���v�
��k{�ɹZ����
C(v��a����k&^����_�ӿ�ʝ�y�f��<�r�p3�p��9NDs�(m�L��x�R��Q5k�v��c��
�;��*d�2Й��]\~ĵ�k�
���QX���߫���3X�O}���UC6m6JW�9U-ĂO���랬���۷o≈Q��L��������>�����?�>����,_���̬�y�w�%��Fm�;��s�~M���,�������{�8ǥ>��pif�f%�)��Z�������@[��L�v��a�55C1�e,��M�5;�H�\���!����=[��<��HƂ2w�u����� S����Vﰐڹ�z�۷�	��oa�8��S�U\)�n��=��� � ƫ��=�Ɩ���%(~����e�����ZW4}������{Z��g��[�ܚҟ�݂�j�iz��J�=ܿ_����湴�4@��9M����Z`��8�=�
� �m+ﯻ��4���(�DN�NBZ$X�v�:e��P9}�5-M����?����nnVZC��j?	�������rPx�kB#Obae.�?�ZGf)7�~����j��zwJ�i���F���V�Y ��̯v7�� .}�"����Y�N.ڢj��YR驧�!��F���x�<�<�⒒Y��]���g�[�����Ӕ�4��	�����t͵����	���]��UX�f4CV-�\��UT\l��-�[r���{YTbm��;�H��{�Bo}}=�y�W�$������Rn�V���@���R	����v�fr�������y��싅|D@�����/B��� `]	�u���
��C��.
�f��WY�P�޿��L�=�A��,�G�y���&(�����"9��b�/\�g�Π=w���'��T�o���l�q8$	M:>^��>W�Q��(��'j�Ѳ���s�t��5UM��y��@�W�,R.��!�?wtt�%�;9!�/H���/��F�����Z��Z���YY��>>>����V*[UC��-�A
�O��4���VbA�����������<����B�=�=�����E�h����ۜ�֦EOOo4�f�!�/�k^�)Q�sl�N�P��)���$�D
ư���*�C#`�`�B��B/~Hַj0ky���ʉc��pG�I'<[��u��R�[G+E�4�[J����M4CR$���,wbb"K���Ȉe�ͩ��U�к$P��;'àҗO>�C��.��fn�
M�����������:��@�`!��t����5Z��$�N�%���׻��D
��͖)�'�.�r�+C�Y�,ʟ��j�v}�[5�?����O{|�����pׇ��A��"��t��_a4��՘��3b�b��3RR�ɀ ���p�v�w��%9H�̝A�M�W�U��ds���G��l�΂�F�%���_/^'*ބ����Ń�v����1+Q�S�9L^�����')���N��w}n~��8I\L��ǡQA\H��
Ph�����^�B򉪹� #���8�,��z�bT<��A�o�en���7���LVq���UB�p��0�,�30�k����A3��鞨��� {�ݥ}��j���-䏐v�t�U��B�a`.���
�TT�1wi���r�%555��r�x \�.9t���� j�m4Ui@��6lQ][�Y�!�s�FV^u&��ҧ͆��E�S<C҅d�f{�,עq�Od�S�gTl�W�?��j����K�0���
�L�t��-�P0�8���stLX	����g������"d�����:��T�5�u� ����a��i֢��o����������NR�1�/��da��~5��˙:ۜ�O�ӈ�_��n݂J��K�î'2G���E���K��"��h8�V�	5�H$���d��}�"V�*."b���? �"53����������G�S؅<�I�=X�in��/,�Z1P�0m�Vڰ[�O����9|������Q��r������`�I�܊���� :*?�K���f��sC�k�+�QW�ڒ�]�����>�гM�7����:����Yۏny�0Y�V\,�%ťfpR�)����� ��O�@�ܦ��3��������
R$��������b�O+T��Ҷ�cA�Ν�]jSv���dC�RTG�Z�$���̂�O~`<���i�b"�H	��Y�����������!� � �ߋ��Qd}����0��i``��+@ϠL׉8LQ@'|��Y,��ݽ��j��u�LZ���% ����ɪ!<�*�Ӎ�%����Gp8�_[��_�.��R�G0	�G�à��H�t�}���&5������S-��оڦ���ؗ���grhӶ#�j��>�����#.h^=��������]��#�����m�"��3��kg�>�����0\���HS������OVy��SaIԆ���9���YT���{���͉qځb<%Ƭ=C'�!����#5�	�����?Y4��Lbecs$Ty͙���7w����'��>��_�<����t�^yE��)�a��������'?�2�]���B�Ho�<؂�,�B��x��,�\�]�����)�J�F�*�6U��1ƕ;����WT��c����r�R��n��Ο� (Q�w�PЦH))��*䋎������s�r+O�/. _�:_�j�v����K�|�W�1��>b�
�qb�$Fw.^± gel�e����/[�\��F���z.&��顗K��;��XE�_����붶��ǡ�j����O�4M-���g�+s�g��#1+3�t�Y�t�/M�T��e��n�����@�:V��ˤ��oYbՏ�IGY�
G����6�'�����(E8(>��z/
&�, �:.>ޚ%D�Jߑ.ߴ�#u
�I/�!v��=�$�/�����"��Q��,�TU?��vX]]-&|���0��,<@�#��H�Ñ����_�'G���27Ot��2<���u�O~���"KrJZ'G_�m>[\Jʖ,y���ޖ�����䱃��1��ƴ��9����?.���c�U3��i��bT�̜��E3x�vF8��arವ܉%R~ܥ��|s���6�!G��߅6�
@�j�\*vo^w�v)�&	_�:$vP��ħ��N���Ҟ�Avvvߩ���?��-�	Pۀ2:� ԉ\3M|�$��NC I���/��sE(���0�_���k�!yD�I!���=�f�����=T�#����o��+*��Dk[h�����ݧ4��ۡ�f[��bç��P�-v������F�	v��k-�eN}�<v����!z����w}u�qF�cSS�QwS���D�smm��V��k#�����-��w#A[�������0N��2PT�T�/���7���k3@���&$��1AY�ĴŦf$�������C<N~�듙���iV�x�����;U�f�T�D$�U�/_���s�[Ip�Փ�*��zu���.by�4B�^2�}����9��<��@9��ě�r䦧�ǈ�6�I���T�OyN�8�KH����8���`��3j:�
��S��r #�F>=xo�]��"jn����ts{MW���%����Gmx =��f(��o������9D���4m>��{!�k��>y�)ƚ�Q��q�W��X�����?���ӝ���g^9HKy}�j�?���\�avW���\�cb�z�h�9�\(�2���ə;���T� �����E@�^�~?��+__I�p$�h�F��y�g��,G8�]p��!�L��k�E��ꑮ7}�97(��j���ŗX�e�c������dVR�e���ҝ:K����yo����׹}r�������%���E1��X�ll��~~4~&8�XzMM`������٩�@)op��
tIJC� �m�l%ZYIu��۷���1v��}���O,=0_{۵eO<.�.t/�+��+ ���A�&�u��D��w���A\�M �Q���7WeC�����Aν/��a@9p�u�^zz�����Mn�ޯz�\'���n�{��.?�i���U���ZP%�rFL�^,�T_W�ef&����X�����L�����}	�}d1		��z�8H��AԶ�K��8K�	i�*�g�p�6_��x?��*lT�s��9��..5$$�af�����K@Zʫ5��,������`
�S+F=�qXY�k��u��������o�m)R)�����7{��U�S�qK�]�;M�6/�j5���ps
op����
{���I������ߜ?y�����ey芠���
��mZ{���x70ٳ���y��l�n���k,!���s�va ���?ѫ8��fh0N+���I (�{�p�=�D��`��H` (̽ T ���zތ�S��쩙_K�=`W�f�}��c7��8������?�����>�4�/^�lb�`ge-�3�{��'%@)��T.�f dy--�$޼�ǉ�bvV�Fc>ie��w2����h~�p�>?�пk]s2`�̬��U+#u��Z-����Zv2�Q�	S[�|8�j�0Gt��WyWGG!o챩e�U�lu��.������'�Ur�-v�#['�ޤ$%�Y�N�]��c���۬3�h�.&�W��_m�j����(u�/�7#S�`(�н��U{�:�Q����i�P&���c�M�ITMh��ɢ�,Zd�ZIQ�Y����ՏN;C��Ҙ�ܨ��k����f��KK��װ���=�9in��0��}O��9���.��BOf	9m����g�L�X��Q��~W���X
X�b��)��RCP
��T/k�^y��P�=����}Pk�6�R,iؑ���>���,p}Ui���, ��G�-�0��Ra�˗/C�q�������iX�RWq�G�}&��T�V��aj�sWɋ����~����;���5��T�$��##�U�ي�Y�'!��d�}Tk��7���g��mȤ���ڮ_`������]�����)������#w5{��3��}o�/~����{��{,`w[d�R�����q�ǒ���H��6�w��%/��犖[N�3����>@���O9�gC؜x�g(x���&�MO�n��PJ؝q�{<xp���$ǡ�A�%�*v�~�Y���ʟ�%�_�0-���36��u�m�7����P�������Hh��h<�_^%��=�6�?=�:8���k�s�hXJJ�7�Q#�׿̲��^���z�Md��Kn�&�������U�������g>��̣����9��e�LLL
���z͚���t���<2�䵸���n�7B�����S�7W:����[/�p�8��Bǆ��oWcH���|��U��}3������νa�9����1��C���Չ&���ש%4�����V�Z���%�����4�M|���\Rc�d��>55�Қ����ݭbĖ�;c�Ɂ|s~�U����Z"�٤�X�o)��ײ�gj(}5��9_�|9��mb��WxfJ6�nk{�6ݎ�-�����;�R��7�afy���o] �Β�~�{4�O>Q�#3�#xz�]�ЋU��n2k�2^'ńu�nߒ��Yo\NQu�[:[Nx1�>�챾��8���)��m{t�� �����L����-)�t���<"�{q�BD��a�s`�N��e�z�w�S>{*b�0�IQ�y��3����슌eԙ��|ك$��y�{Jȭ�-,��s~w]��Q���,6n�؛��Y�jU3�[�M~�.ذ�tBK+�^���iwq��oqxUD�q����^.jwz��u����D}�}3(HM��x?%Ȕ����$�0Qf�T�6�{N�:5oH4H�)��{�.<8Lt`g*�i�,1�3�z�J��Wџ������G������.��=��OL2�<M+�ߘWP����d�?��!gZ�w_�~��t��T�-+d�����]9{�) ]�R\�0�.=?�X��E�j��Yma�ۑ��	����j|"�����F�_e���Lkb�8���1� �x�R����ڸ���-�T6���+�^�u����!�ܹ�޵�����v!%��#�K�o��/�o�&�� GRA�~ҿ��[;�[�����
�
�L0���d~��Uua����`S{{�6�2�-����6��l	��;`�f`J9d��}C�;J��&�F�`b�@���K"�5�v�p��%y��]��-�XU__�e�v����1��ͫ�-o�;��6�.f�� 0a�#O�t��u�U��X[���h�.�#OD5x���#i���Tt=l�+^���5k��G��R�a����h���<첷ظ�,�C,��>�A���0�����v�v�S����Rm������UKˤ�"N��knRo�*���l�K�y�(����s��f�x���4�z.A�
��`�2�G��Eq��o�vuu]6�Lw*a#�%��k�w���E������gu<f�Aa��-AMCÙS��\;^�Sp�z�8W5h���36�M����5\� �%��6gT�D[���Feaᘻ��^�`��yӏo�Ὓ�v>���{��8g�7SO����@�V,���%�W~x�^FFF{������cfڔ9�@p��������UEE±g�D�.������Ӻk��[�f@\;{���p9��8潘m������+��H���A$`���lvt��/�ޏ޸9)3������q��Ys�zZ1�t8��#���3�~}��DeIߒSr7y�Iug�����eS7�7��w���B��D�k�������"5p�ܚ{!��W�Wj8mZ�	z�I:���'��5Rr)Us�ί-6�il
�w�t�e[ll�ݻ����o,4�I�r�3�G�|Ōs�31U1��� ����9]ōM�3#3��/x��.'˳�]�>��]�)�iF9�n���[�x|`W8f�rI_����{��9-#��&�h.q�/[���B+������)�R�����Cr��OE��k�'�]_�����״���4��>Vn�Ft�m��V�E�7~������6sw�&���H:��{� ��}��ț���H*���˗��k�(�6j@��n���y���Q����*���uE�%�z��3�f�?����־���3T��ᗽ$^b�) _s莗�D�l��y�t-��B#�
�ے���ծ���t���y� �ے���'ܷy擺ES,�����rF��Kۅ�!�m���9gzI��Clll�_Q<�Wg�j���ӛ�.�<0P=���u�]��r���a���Sp��1]���Z�Кڔ���Z��۴�߶����Zt�)G?����W�����"�Y�������z�
cQ3��%�)j$�}�בz�5��5� �H��(�N(�����������Bss3x֩$��V*i���U��<CԦ����������xR��i�˱g����홗ް{� ��$Mg��ɔ���υpǜ�z�z������Z�`��|���L���!š��!���u(޹L�4F���c�.ԗ�ڈ}�ė ���W�d�����([�_�zs�_�)8l.p���WQZʲ����nhb�~����������{6����� ��n������h�c?SP#m3��\�K>��� S���S�[Z�;:t�y���t4����D ^�oi
ۧ���<�f<���i�[g�6c�J՜��&9:���S�_ꢍK�&�[���ϊ�>�Ȯ�_S��4�Rc5 4�Ibb�^H������}3�2P'T������	~�A�j�Ο\�s�h!D�R=#e�S<�?�7�OU�aF�R�54��2&�7l�׼ߡӟxs��a3��#� ��^XH��!�2����qo_ѥ�Q�sJ#0����������C��?��S�5�j�G�$�?��y���H;�0�@U5�Ø�Q�D1"��V��	i��P	��5���Bϡ���B�5k�7�;2N�����֋�S�@��R��{�>�8_�����Σ?��>D/����79�^�&��x��Q��ov����ѱ��K]f0����;z���ޑH���<�J@��~
#c�VM�.$����jl����6�rU���NÃ:U�Y�n�%�[>}��U�b�T�N������,��!�5���%�������]���v�'���<�^UXK���j5��� �ba}v�:%n�@�z|��'Q�X"Ba�����`jj�k׸��
��@Cw�Z�D��,�/�7d����(���/�����V>�������T�޷"�� g�^����9������3��7!�����9
��6����5���gm�@�=�_��_�L%R��4v�#ú��F�v� �ɚ�Hm�s6�A�-�q��|������1G#Χ�/�����fo@���Qs�
�V�E��`N�C�4.Ҵ�Rr������l�R�Yl./,�5x�}l��Q�	�&䣚δ�F��X���T���É��A��U+ğ��?C�6�0Q�Y"S��W'#sc�c�"����w�ȸQ�%ǻ�c*��ǈ������"������Γ�7���#���"�~�x>�[gv��o�ҍ{f!��7d���!/$k��Kg �k�4⨮炔�z�Ib�"He�?�;5�(
�\�b@{\|۾�0����VN��mtp�p�+�0f�X�F�B$Kxå�#�R���54 7.�����(i����R�a��v7q���N�7�3�	'��ܿ�3���mvd:����F���bu��km)�ڜ�/�"I����:�JUA��<"�n����EE����Kg>~��Ms�H��m_�IS�R�N�����[Zb�Z���kn%���)b�f���-���w����^���h��J�³j[
�e�vG$ԏKgd7�/u�� i��/6:�w=+r�Ntέ$����-��VƈF�P �����#�s�攳:/Ǎt�q�F�Zy4� m�{����{�X�B����U�G9!�R�8��A����Lx�FoT.������J����B`v�~SF�$�2�0�
�����>�N�iص'淹�;�?�=<�$��/%�8�^�5���p�l�!��N��"i�)"��[(�R�F����1<0�p�I�#�!F�D�s��j[q�U��l@��U�S���e}���zT=��x��R�W&
i��l��d�c!��l��H��ٽ7�
�����n|�QPa���m^A�M��~s,�K�>d�E��G.�QُC�&����h��Q�.{ǎ�����z�x~�#xx�EGY����� �iϊ�����\\@#"�͖�>8ȸ�������<�����}1�j�5��C��،��`�X��v��Qڲ�J`X!�����{����T*R�m�I*7�iT����鷟>����'7���ݒٷ��Ș�e֣1l�&�6[�;u#�!�s��n��)�灆EGG�����~���Kx�o��6N��ߒ��mBڿ�g�M��T�_:>>��3V�Y�i�*4kԱ_b\�r
����m?T����;��L�@j��!26]�2�E���O�Q�B�8b<��vl�J�|A�u�՗{�X�u���:�rG�{ն��*��c�&�H���ze\uh�q����/������06b�1}����<�3��8S�p[�mx00���D� 0���E��;���\��bbt�7�KSs�Xl�ۥ��?\���� MM��-����&9���.�m�
�i��/���҃+����Prl������NE�ݳ�]~W�i���`�fGN���]*�%�Ner1���J�xK�X/�{���t��q�g���g�6�VoYuvK6I�߿q!��ͦrR��?�����'rKF��!�2F����5N��s���<Z�N^��/�<2�G�.X���P���˙��Vǵ�K��Ϗ�Ќ븄�`Ѡ,i%���f΁� ��,6��R��W&�Ŕ�E�����&'�-*^��*U.�/���G�H��:z:c�����v�F��r��R�M�v�N�����w����Db�� :��su R�ơ�'�K��E��Iu����,�~�P&��-�X�o�<�&h��&�;]+���u�H��<��e|�8Ƴ���$N* �s���j9�~����M��y�{ґ�_�����_.Y�O��O��1�ׁ�M����?�m�y��t<�)tڍ l?�X6�P6۽i��e�#�o�)3!�W��a��V�M�D��)Rq��ڟj\6-�?�V��L}��dϤo(rt.3�������:���ЯM;��p�������9����`Wd��at�X����;&4�-�Lj*;�h�}�;����O�_�6�h|�b��W���`�����Դ4eoS�!jb�"�ɟfs>Up����[�SV��@n���2�8���(�^�o�3g�@a��t��u4D^�Y?�O	Ϗ� ��RzD�~n�f)��W&��ƪ����Ǻ{�Z�DCQY�����GE$#��]���<���d����P��d'�{�����>���}^�筗�=��u��{�s�<س&s�z@�q�`AO�/�:����#����ƾ1l��une璻c��+jv��ݹv��{�ǖ:�I�Tc�"���{��.�k�*G*G*6Fn̸���(f��G����4�1@��I?�kT����uZ	|-0'��9�m|�a��ᢦ�|�#r�#�"C-�D��3�0Y4��`��J����\�g�z<\uw���%����M���W��ܙެ&�p����9�ğ1^+/2��b�]�����&�br���m t>�C /n��a��t����釂��W�sH1��mee�����k������"k�b��&��BL)I�'��k��b��Yhц�o'�b"����\������qhB�J��a@�XBn�j�T�J񄔮u�����/$�޺���(����"�pL�/�Vi�$"obգL&������70�c9o?E�t<��D��{y�-�_2B�+A��4*	�M5!U��U�����jf���/Rc�A1Ld�"X"|��#���~5�c��u"=!�O(����]���}��\T�
��N$q^&��E�%�
#���\̨2��C�1u�NJ�{�n�d�.��^�@����}%�g�^��~&� !�;V�bG�0LѻW�C�KHSj������~ʯ,orA)��0��þ�$���	�B;��N�G�~'��d�aL{�Hq�ڹ,���P�+�j�j.��R���?�;.&���RІ���۷yLg��U(5�*n������3��':��
a�ݸt�3�Ԟd�&�#�b�E>���e����v�B!`�%(�r/���r�3;�nr���c��$!�:p?ӗF~�=>>���U�)�`��I��~������w-����}9pᗡ��:��EMo���'3*N�=A����� ��"�s��&��r��h�'$�Ø1�V�	�ʄJP��ޚ���'(�+o�1P���pc㕦*?�m���X}[����| v�O��&�Ҿ^���^�Y�t\nb-xlw�p�����􍳩=�ō�V������	J��Q����U�<H���,*�`�2���}�>�&<�:/8�Q`��s܂�z%o�N��R�b��ЫD���7�a<���g���#���bf�����|:�����YEL.��(��~��,��fΓ=�.�b���Ƌ�����)	n��M�(�HŠ�ld?5�bl}cl�!שR$���}�Н�^��Nn�[+!��LxZ}_�~�U��U�]'Q�ƣ'�]QϢuP||S����p�)�)(y��(x_�- 3�n9�y;b�s��0������G��*䑆�4��\��y��\�_�xlv߉p̣�bc���ӧ+���y̤#��(���3	�oҫV7�׸�[ösnQ�b���֭�YY�LŠ�1�KX�8~���,����Ezkn���_Z��O�/��3�(���z\C;��ܱ0�sI�#E�	��V�wh�B9��?&��tP0�?�	yL��ɉ&6�Z3�lrV�����W��e$�>�*�sg?������پ脱�#G6��u��e${IV�֐�3��i|��Ȫ�n���;%Lv�h\�=2���{�i~�$����=��T�[q=�J9JW��:,r)�˹���:�&EF	vs���Osw�\�mK~�d�On0T)�<�%���0<6O���c�� f*I���mL{+&������S�LcI?������	jq�nQ�%��#�l���]�d����ܘ�UX�u�}�����;
�O�n�QN[����?7U1�T��D0ڨUp0�Q�P`�S�ۛo2�{,МH;����ų���I�6�Ԅ�X���]k�����I�	$x�|%}�ki�d� &{/Su'P�ѯ�+_-˶�B�����r)ʁ�$9w*��c򟝜h���J��)��-����ZL.7�j��5.6���zJƝ��|��9)��	�D�O�XV��vb����'�YZ�Qn�A3��GOL���^J	?�m��y���ى%�k����B����Ŷ�'�ʛL[�nَ%�Yc\���k�$�N�C��En�oR��'���6���4��F��xWP
���x*�RMY�5Q�w))!ۦ�|��V���*�cOp$�[{go�N@�M{�O�؎�ib��W�Dj9�wG�1b=/qs�;�u(���\�~����GOH�8�t�?��QI�- k}��D��Tl�$�kMM)��W���7�`ҟak�ZR��[	��qf�����4`������X�6����t��~������H����f����j%н�=ֽ�l���}�8Ĳ���O��!���m-���*�����(Xz}L���!��ర�RK0���l�R��_ܪ�Qq�LPW�}n6r*o�+���g`����>�m�`�iI;V��|�>��.��S��66�O����+�^���]��e������p�-�m�	������lł���0���(����$� TE<ҜM�S��c��n��x���%.$��ؕ}l�È#��mD�ƆômO❰
���hZ���jٳ�9&}WD��B����{m�����HF�?l_�_p�'��ݓ��x�����{|d�֋��Qу��n������t?V�Qa� __�@;K�q��[�K8���΢��ע�)���A�j�� ڮ���z;!8*�9�͔��	�t�z��S[>l�ā��tO&��:�j�F�OW����N��Z�u�E�싷
{�Q��� V5���m7Wc��<�n�Q�o$�����������ژ�нIu1*.ȋ0 ���b�S�����B����Ln��<̟�s�C¸�lCG�I�ku�洴����b �p�&����]� �R��H�:o��:�mM��?G���P�:C[6`������\�V0�)��BC]]����W0�`2��p%��b6�L%��
U7尛k�G��X#�݇n5�WP�]�^��Oe��hW1�TQ������ŋ�*���ϻ6p����Og�h�]�jZО�(��{��^��nQ{$�<}�RKӜ��8��-~�Hs%@�" �؀ln~��_�i�NUUn��O#蔖�q�E���\Ksc����������R;��1�\��zaL��yN�\��T:�}�^F���Ke0L��qs}8�xgC�R���x+�Q�>�޼M>X��^���ܖ��Ϲ��bA%�mP�	���R�����kZ��>��r�EtB�%�cS��łI�k隉��}u������s������4.J��!5zj�mjҚ8FXoʯ�?_8{���BI�rd�}�e�눛��֒���5�,� ��~7ġ�p���'B#E�ï�H
%�N)7{sd�t�!~҄�mNcT�d�ׇ���r�⪪�ህ��0���N�������'�m��S���檻0Ҡ� �1�_e��@	���6�~@]�'���`�/�����[v�~OJN6��n���m��������U��Q����K�t�ä��g՞��,��>ϡ�[�ՙ�+�)��u��Zƛ�!�>���

����0�#rl�O'�%6=��k-��ln1D��wߏ�����^�Ȥ�n6GV�0.D���k�g��d�f%�kn6����|�A����;x~��BT����+��f���Y��z�x��k�G�̎�w�n+��ɰ��-Mr�ΐ^�u��VcDA�����/Z�2�A�Ң�_�SGL{엚rz�f�����5ʽ��lOz�^�R������묯����w��yf���;�.�} I>���۳����-,,��Dh�/4�o�#t�7|t�H<�j��O	[��fZ�..��btX�j�d��9G�i�����ӿ=�j�[���)�������W���6�ʷ7H<3RSSWF g[[[%^�w�B(u�H�et3a
����ʛo�x-�`�ky�i��E,��xE�UsyqR��X����.��t��ǭ�x-�nt�fK *6�j� ��CFgg�>q�����_��*���'1��{<���κS��8.��RZx)H� m
��Uf��^��H\�z�|�n^RW5���Cp��A�����,�1^rn�����o=�v\���<��Oe����dCL��U�|��N���c��D�BA�����Y�[��A�V�Bڷ����������_�Hf�ɜ��M�b�BHn��oq������9��`Ŝ���QF��y2��3=�~�3��z�,��$�s��w���I]�l��22<,_�X�˥ߨ�Ǩp�z2���VKCg�����.¡|��s���c��y�I,�8:F����u�(iX���2�2=���CH3�M� k
߈��kj��EU9R`��='y�����P��e���Q������S��C"�÷pm��"��)��^�E��XÈL����xY{&�z(��/�@�r�ѢH���C׽GQ燙���yi瀋�֬Aq��9��e���<�}@�i}�>�[�ī��� ������de�MjK3�N ���P�7��P���`��U��x���N�_�UD��jj����������Ϝ/��	7j�G^���.�2,b�2�d�kPlJolL���mL�����ws>v
b0gz~I#K@�ҋ-j���nQ/<=�[f]��t��)e#tF��r�|9�1i7_�Y\�=0�aDm�p�Ս��M�NT�k�E+��-�x���t�{�/}���������B��':�,i�LqQ��G�H���h�2��� �;H�8L�J��
8���{Lb�������}�\ٝݍ-'~r���z��◚�X/��1o���F�ψ{}^�磍�����!�I����cű
&��?=A-�7��X��x!����)���Y�ېfA���D푙?i�;����;!��Jm�
9�jҊv{�lA��bjtp߂�xC9��kW�lG���K}�d�H��Ԃ� �9��ѣ���	�܇e�,�t����F'K-��22�ҟ]W����>��0ʕ�)�M���B_>�B���lÈ��������%���e�a����N�.��:���𝞼�W�|�[��xRfY�e��_�b �s�z���|�D�gk�	���Ap��]���Bu�����|חEC`K�Ս͌Z�����;�jq�hq�z$�*�4fZ�G�2�2ii�Ŋ����#/�\&͝58/^<���|y/_�W���m8�eG8u������,��kY�2:�(My���4��v�$͸{�������-`�T�u�/�\юl� �}@�az	��������xr.+�ȡo[2U����}R���A��!D&�!z^�Oܛʓ�ʊ���q�̐Ʃ���'����7�wVc�5�y\�m|��V�Q�i e��/Pj��x������t���C7ϡ%�O�;����Q��!�kb��a��+���mo�F�7\~JF� �U�=I�_���/�&���A�����`��?\6޼O�o���u�ten�Ҏ �+����]��`���.Z|�/b]{���э�]�K�~��i�_��o��51��*��>�6�O��q&��L��>T �a����HP�sB�������]v�s�ϟÚS�'-�;�'U�:F�I*�����~������z�B\����J�ka[����!�[��D-�Ȅ }�l����{r\�7[u���Ð�!�q)Nx�|*'9Q�8n#���%$�_k�#�5�~�"(FE�\n:�(}s�s�!3t�1^뽘�)J�ii��Z��9Q��*FX(:��,��x��2�	22�򊯺\f��_Q��0Y�P�2|���-<��R6�S 2b��֊�|U��V�2��2��%�*p�Ĳ�afǢ��� ���CCC���5��Q~�)%�u��tL^��<���x�`6 %�k+�-�,-͕�jLx�x<%O{�w?��G�$��7�����T�R�ٛ�t�Q5�,S�uKV��i��bJ��Q�6E ����� ��m���B'Pn��)��3H���@@�>|��׶Y�.���^����گ�{MkX�=�{�w,ɛ��	�ex|�zy6�DA3٧m4�R0��F���FohJ�Jjƶ���ӟ!��������ߗ|����0��->+hH����)��8�k�KY+��0J�d��3>���O�t%��j?C�"�7m?}�򌁟_�\�րә7�Vj��������T�k��>x~7���Nx��0R��.���Ӊ��ۅJ��/} wtToK<`?�a���Ą״�m:����yMW�Ź� ���������9#~����ڴ7R��c)�����\�垐5�Q���Y��LNJ��ح$;�/�>Ik�� c	���F2��������C��l�lٹ��~-�G�Vx�Ix{M�^��s\�_��r�U���66|�Ϋ������}�:����dLC�igZn	)�N�2�s�������)��4��e0�d���6;�k�_����0����!��k�F���1��k���H�����R�N��f�


�����K�[K����
�s��˟�
`��<��m
�a^�j�PҠ3��~�t��ŋ�*��� h�Z�����Ͳ�z�AB�CP�� �=�т%+S����-3xN���l~�X6\ ���x�Y���6�I0�La�7��Db�;�k�W�zVYlw*����33�رU��H0t)-��s��|���2�Tx����詐� ���7�r��Ӿ��Y�1���~�eo˰���!���|�d-�څ4Y蝑��/�JÉ��\VV��xS�m���4�D�~�Dm��>��n�#3_8k�C�."X ��A��erq�ˬ�e�׉$�KN���۸o�1UY:[���5��~M��;O�������M�ƻ���=j7�

��{0�o�~!�-,I��"G*ʇ�/_��:�`"�kA��CJ�!d��?�15�i��@yTw~NJJ╫:-C7���~Bk&�Ğ����4�g�(�d�OOg��ED��V���4�Ʌ�)_�`� Θ�dm�m���GǙW���T�����2�MH�H������9����7G�7p�%���B������ƛH�0�eZ����*>���[nl>'�`�=0��39"����StE�Ϭۢ�SC��&�V�;��+:K��^��sb���mug���,-HK�k_T6�jA^n.{o�R~ ���khی}n�B�˴���,�"}�>�f ������>/��N0���R�cM�����c��n���qcY�яQ�G������4����]|�>i5�^�;Ӏ�z��q8���&�:�i<1� �㼸�?ߵIƋ�Ĕ�g	�)^8n�l���^-�Y��Y��#O7�I3��{أ��ivc}�x�b�<�5H���e�2d��+3�>�2�i<�@]��Xx*�_��ml�	9��m�-�$9�� _�׽5�����i��[L�MM�7�
�,��'�8��򉗻�J`qkE(4����d�Ӄ���v�w��S�=�6c�/��5�m��b��2;<�Fj�J|0]v��V�~�w���Z4�6d�T:�E.^ϼ��]F-����3ގB�u�q��V���#��駪q�HI+~�~�R���а�k�~p�~����qO�!ćЇ/�=��&.��̓9Ξu���#Z XS�аF����Z2z�9T��[[_�T�۽ F�2����3�OyR���ػ�zYd[o�9@����%o���r��z��oj�:?
�O��3���A�k����y��K��^c��q�3ޔfff���u&�����ze���/��8����F�0�wIIb)-k[m�s��S��s�]��\x=��?y�!�̵���D��2����?{M~��΁Q��2�<�ldhh���|�P:�aK�kF�Ǔ"4>���)�;��Jp��kM\��B�U8n�:|)эibjs��dz8��jG�qAw�M-Z���a|t��6�s���i��|�������2{b�Y>ټ�n����fJs�l<es,%�~�)���q���=܆_ѝW�)��;���x�������
��{�����ɺ�󩏭Oݣ��+;�՞�ͥ�ر[��;D�ƫ��o3G(�	�T�AAA&FƬь��KBڻJ�PÑĴ��QF둲��tQ���K%���T#q5w�Y�f��L���`֜���$հ��&�����k)�S�˵w�5��)���D����Z��U'���4��y�����19%���$�<☼�˚yzo&�yϐ���o���P�~�}��r|�����"�6P�]�*#{%�ޢ�Y��)=���#.�������=+^�l�2��Y����U�9J�Ϙu�A(�h`��:�1� Ռ�u��X>|�6�cF��_}�%w�����,h�� �g��oSS9������%��!ܑ!�r��KI^M7��������)�i�H�5��Y7:nv<~(ZL���¾}����[Zp7��D_�=nue�9���ɀ4>��c:p>W#k�Zm�,(5��3��.ԙ}fE���P�[���ʁu�^:ʒtGv
#R2�����6<6w�l��@��;l���Dl�L�eF��G3U�HO�8��Z	�Y�}���ų�	��8=���K[ߠ�k2�&�s�jVϵ���m���E��˗�����u�R��N��C]'�,��CQU��%S	��a;�� �W`:^��L:ka��+��s�!!-�h~��Ӛ�'|�L�5��l48l�?�Q�U��j��yuę�&�>�Ȣ:lN�YV!R����7~u������n#���{��xg�����Օ$Ag�|����Rfo$��AKr��7�qR�lmm����@=��-�`m���?��#Og?q-���d2ߨԖ�p{bu<͈yyd��������mJ�������׺lzi<@I����B��SS���BK�K���Di}9���VH�������	�W��؃�Q��`�%sai�����=xܳ+v�T�
�L��b��ل簐��E���|���,��X���@��j�N%�4����t���sթ�;�'�n汯UԨP)1���h-��}<���{]N���qn������2����K���~-�����f���egV�W��$Y=Җ�������\��� �(�����Dt�ي�=����Ys�!�	�����,��Ũ S,Nu�6�h�>�B���)-y|���{e�FG_��JF���G'i�Ěy��ԌU�����k��3Yu_�J{�;C�&�t��C�';pPF��B������h�i�ō��y~m��#��=���ڑ3�$�W�وP#σd��|�e��Cՙ��Kk���t��]NO��d���d8���p=�J�$�ϵne�}��]m��6jN���}��l~MY�=�Q���P���˼���E}aǓ2!:��O�s��ͻ��ʠj�@&�+�~(����9��Kd�
Y�$�F�Q69QBJ�'=B>���q2ac�Y��)s��}|��!��>'��O��"L�ê��[�c�G�m���S���3��Ůk,���T&�4� �gÄQWxz}��l6�׼�����h�^(d��(�h���W�l��裻2;$#��g�@
��c	���N����9�*�l�� ��)�{�:���p�O�I#�t�����,,C���<@�����g�W\��A�)?�|I�2op���k k���Բ|�T�M��|Mx��"}�=̈(�2�aW�x�������+��8�o��s�!N�5�|��(.�����5����n���m�Xc�\�pHOK�f=�s��cNn���{�u		��J�n�-,MuA���|#q��'I�c�(#�K�/���z&���ߪ/2GԎ����Ĉ�n��I���J�vG]?�d.!H8�c�lhoo�����I'�� �^�#��1���i/��m`�kYj��	��p�&yg!!��Xb�~��}2��{_ǡ+�{�r���p��W�n���FP-?jF���Ĝ� �]~ɨ�;̓u	]{ak�B�߱},�z�>��������edn�`&"������ U�EG�qb�_
�9GJ�#��s=e�F��ÊN�j�W4����б�5�#Vr" �7#0Q�k����w���l����цh���cc��lO[Ϛ,�5�z947Ɣ����V�K����0��ʳ��"*o����ܠC���/��[���
�1;��=�i"�u|rCs�1<<L{9����HC}�0��E�Tv?.�$�?Oy�o3�+n�[����ț�i{�m2 n��Y7����p�㛜 �z~#��3gc�)��餤��9&�z��t�:ZR�V����G�3�]��;:SN�R`��^t��������s�	�Y]�)-�nnnD�C!��:�113S`�5:|OWUU�;ƞ���)�0�I&Ӵ��"�~�g��d�bPm4�0|<.�]c�C�CS}=ǘЇ�w��ȓ!�3�[9a+��ؓ/X|����=���6���$������s��M--#�x'QCta7��O�K���ΑkS��ODD.^�(S���2��8�НoH���*}�>�3�X4�	��kϠ<��J��h���+�<�Y�[o�d��'A�Ae^���8住��mt������n����)r ��D36��CXJ�%�ȹ���M(L�`: �OJ���~�?{m�gOc#��//,.�g<R�L���Z�^��j���'�cA��m������Ջ��P___��56(�(vW�xNU��١�͖�sS���F(�.wO�'�B����7����3�<�4$,3����OЍ���i���� �����fV�r�f�9�5%���2�A��T�&Y-�e�h�ވ�r?wb���F;b
�޿Ő���BMt���=�qYY�х�i�*@ƥ�N��Qn~��큨P��Z��ˢ���qRҘI
��G�_ �##�c���7���W`���4��W�$�x��#���f|n��˪�J8]��h���J�v�(C|^�ڶ��jг�y�����B�d��v��
G�N�T��}��ζ[I5Rz�]z/�n����
 �s�c����}4�������d��g��-�A���������rv��U�;
Տ��A��9�����[Ǻ��}�k�%�����x�5v��7�ᚐ��A�����+&����L�<JByͣ�@����C��	j��眢�0�#~l���#�z ����)�����n1q[��H��E���u|r��c��Vp����G"�+q׷�k��:(��A6,Tkn�ύ�Z�mx�����ш4�H'rHt�����9�@��f2֞_��t`��nw�ˁ)� )�LL���mo׈HH�������N�k��?Yq4�۸������(B|�n)O�iJ�vqBE�>̽Ш [9p��4xA��r�횕 �C�&��O`�����N�5��H1�w] ]ݝg�Atf򵏵��b�x-r�c��vŽ�N ɁG�`�; 
$yDhހ9�)	���7�|:h�����r���k�=E�]�QR
Z ��S�o���Y7���Fq�ģ厓��X��*���Z�is�;;���@lR
X�\[��﯊H�I�y%}d>�Ň��{�sOr������3COOLJ°���T��`<�+譣\w�q>EO��L^���G�g��㣢���3��!D3��&�l�/N�q3��=��*�6�47����?��{�Y�Q�ڔ����|PÇqt��N��@�5uu�wl��d>}Y>P�v�9CV	�D~�y8��̰~��8���/�99�	e��t}��w�#�D/q!1h~���3Bo��$�P�Hlll��M��}� 2P�1����m�(�gGF]ݾ#~ثAV�u��Vrŏ?�||�v �%��oT�Gm���߮:tHoq��p��8��b�����uu}�4��YH���u�d�+j�>;k��`*3N�Ԗ���uX.�3�\&*1�#�x����x:�n�������|���9cV	�1vB=�J�8TL�b ���3�A�@�ڽ���-�WA�� Y���wo�J��˨]���_�l�TR�]�h�			�D��my�s��$*�X�rНp��L�3V:-�l��2(��_��*���q���رN�x��P#DD��\	�>]�~�A�����-�lH2���+@ѝ�w陵�[��oe+����7FV��|�1ð����]x8�9�A�%����x�}��0�iq������0����9�P�����ysG�t�ɓ]5z�V�}��QL��
`�g�/j����Ȕu!��y���I)Ǐ�C}�XX�V�Ft�|�ʩ��C�Cz���"L}.���f/�������3V���թ�W#�m������J��b�s�D1�m(	��K�R�� �	��3�,�q�cc���F��hkBy�?��� �ş�y\f������w�sǓs�?FlHA՞	�z7N5B��N�R�C�$�rJ?b� ު=)�nrz�Z':c�Z�gW����J�\�.--=)��[9��J/w��w���(��#�X�i�_~GP�+!����X].�����Ж�'{ж���5��-�Kk���[�kZL�p�:�N}&ˎ�ˮO:��+�<�EFJZ���Q����S�*�	�.�%RT_�*�I�}��!w�ڣ�E�lu1�0I��4��c�DC�JX�Hu �2�SˠR]h7HA�����ͻ���|��c��O޺��q��-%qb��O��JG��҉E�ռ��X�����k8���^�#{+&�Į�� ����J� -�ڮ�̟?s�C1�5@��������y��
�K�Haa�z�J��k��:�{�٢��^(5
Vx�����fӄg�����)�c	1�>1Z�Oع��@��М��\BWƂN�:�ݑ����t�ܹ:�gJ����9 ¿�������r�(�u�s�=���Fe5:.Q=2�KI@����R˫�|XC{GGC��旕��tGWz(�u�<��(<��b`�'0���RP��sG���C6X��g��S��H��9�_���NH��N����L�WP���q����OM�Ał1�P��!]�9]V�2�+�u5�G"�\T���(J�U���妉KbVl/��h�v�Kv	?i��/"Ym�*�]%��N
��!�0*��L�lD�UbT<�������'�QS"�����-6rs������WD�Ń�cM	�_ �PbO��0#C���^O�b�6��ţ��^�xFO�3����N-�Qn=�in��$*z����ĉ���/3h+!X�|=�$�sdW��8�/���_��D����z-��P���Ꚙ�f�����@0��4=��'7����~��Hj�F��R�A�������ht�V�(E��X|�G����m4ᮭ��3񮯗�n� ~1t�U4�koL�#�mV�6\pvmJ�?S�~��eٓ��Q@A�U_�F��A��_�d#)�Z��k��p��=�4�1 �9|���F������+xy�̶`34��zD�&_�~�]ܯ��|%t��NJ8?�C�|�E%F�v�-0 ��S=�4!�AA�V��C���l���abFX��\�^yCT�u�ۻu ���c!~��������|��mj�|�C�m��-��=˴��d}��֎<+��0D��]Kj���2�B9-����G�D1Y-�����իW��|Gِ�P������Ru|�z�H:�rZ(V��nQ�¨�� �¥��yVr@PZ�-�c�Kݏj�O�_,�q|�G�Ca���r�/��@I*���]��6+��F���L�5B|�K�[����5���Ͱ�y��4��j�`���W3�ޯF��y���y�/num��)<���ϯ~���	wu�򁭔����Dd`+@�o�.܀���`I[�޲�5R+��Ԧ9�*gm��P�����X�>��Q��W�T�%��A�9*�v�A���Qů_e��y(�+a3��X/����?�r�I��*I�����0���;��e��+������K�%y�n�w�ܓ�=��S��wLLL��6�+%7B���jv�4�4_�1v���2�Iq�C�(�ت՞e��h�SN((�(����:nN�I��0�0i�
Hj�G�Z��h������Fm�pJ``���Sg;2�����7_ؾߑ�2�ٖ7B�#sz[��`���'����(�ee��ra�º��� ���G���-)ö��-�Jc�~ �ՅǤ��k �[��sef�2+��6s�<ljj�v�N�1�c�[~�M����dy�%+�`���/	��4��z�iM�V,��q��ͮ��~��U>O�5C��V�m|���|����=�?��19�s�ZrTRP��Sޜ���N�6��T�z=e�x��F���|�/
�(	����~R�Ь�g���:<��F��wxTwJS�����ש���$�n+�(~���ӍP?�c��&�Bi�����-��#�	����<Ǡ�趝Fr(b7@S�s��T�N���QV��J�6�&�(���d3�b����d���\}�S(R����9ȜR�O	�5�[ݘvLinV�qœԲ�Qw5�C�լ��(|���& �M�9 1`�������ث@%�v���؇7��7�g���.��;�U���cĜ%pC�]�'ʽ�b'644�ՍZb@�����4�g4�#ٙ�W�t�>A���^����w�%�?�Z�շnbK�N����HK�dy�Z��������Eս��cAq�
�}K�;+vB.Ǻ��������!렞�Ki	)�UA��²ZB��FVhE4N���@�9�ҟ��\ʲ�F�qQ�STT(���S���t�+W	ԯL����.%|0������ORQ5����#u%u/��+ U``22�����_�����xG�rJ-I�#�g����������8B�Io��@���.�����EGІ�����8hN�z������N�<�]��� /�k�(�#o�~)_���#q4Y�k��#J{|C ��m��K����h�
=��z��� @ę���ܺ��z�GbV�m͕*%d�i����|{{�|�����h)l���'T��m�lB蕇
;j�������]��)�ո߉C�x���ʞ��6�H�h�:��f�4��v�և.T��ӓr��7__6E�٦@b�T�ʣ�mŗz			C����$��h7Oܛ
"��a��Q��+t�b�;_5��˖q`R�����˰R��u�����d�\���s|������\����������O��Dh|ʴ+d���Q�OJ����+��29è+���q�?��9�L�`yf`lr��q��%=r?za���F�����f@@ P�C�g�N�M)�K�����/E�x�k`F��䌇��,��4 bk�p��ݛ�S��#*�v|	��b�����j�ƛ�T>�{N�D=�d�7���ߤvX�V�r"Uy�	Z�ǜ�$'�����ӥ3��J����c�XI���k6ڠ!$��z��Ot*�>;.���`��3�̄�@�C:����@�t)Z�^���
���'���!��q�U"E,�I��� Hх-��|�v��]4����\_�����|'vj���6s�פ'�R�-_RR���4�����`>�~�?�4�]�v���x`��."/	��	��� @��"R>�� ����F�Q_�f�FuЅ��qڿ�Y�#����w�F -���&�9II���鹌�����$��xy��̊�̀'��]�?Sz�L֧���LV���ɳ�Om���Lsr-AI�N��Q>P(�e؞~-�KL��)��T��pA�)�4X`��[R�@
A	��–��OQG'6!1Q�0ܤ쎝�_҇���JJJ�z=hioOpvv6��"wNHH �w+�l��@C�C:�Nww����RHq9�,�q_c]�^ZK����0��q6����4�O�Z֛��Km���B���G�'ڜ� ����/w��5��$&$�fs��:�2�UH��'�n�B5S����QuM͈m�C��"l*�n����M�ލx��ɢW�WI���<����Wkn��;8��u�ڃ=;>�:}�@ثءm�H��ڔ����sz��r%�@�R� �B���C�bo�U�d����K��N&%|~KNu�L �:l��<����c�_f��䱛�;̔�RPW�W�V7�>�_H�M�^Bv�2�s(�PO���܏SN*�,�ߋXv[���T�?�g�_A�y78NEE��۷7  .^���Õ��N��;�N��.l�:�1Z,�aʃYIPŀ6��5���B~oSR.HW�?011�D鞦�Ǥ	pi'�+������gY_"�5�Rd���䃨����Ea���G|*eRB��X���B�(�Z�M��`�_G���D��=x��L��	9��6P���^%ˤo�᳄-/�!r��Tt�� 64Y-;
ʱ��06m�A���}�e	v��1i5��ߢ������`�b�'b�;�c�9 x(�����t���!�<� 8�v�ѡ0D� ��Ы��$"�k�_2���>;T=����w'�*�i��1y��l�ϡ�������74��#c���J�;���:0֔8 �5�9e8DO���'��ْ�a�\:t���7�C�|��R�/�@e$�<q�壘��}UZ]V����"WL_�]P���..g��
5uttZ�~Z���Flfs�7��E^E��2���/Cf�OK�/-��~��;Z��q�5d��;j9EE�����~���_%���A%
L�d*!k\��U�{J>VS�J���jEb>v��3���j��0EԎ܌�����pVf
��*���Y��ݩ�<�߾}[ Q�*2N�*�Y���uy�k�5@� a�J� �H���&/[8�����/[O����aWQ.(Z��Q�?�Y�%��h[�r���oz��h��'#���"$�����UODzmģ������,m���B�/��|�D��|��Ѝ�b��/7s�ߧ
~)o��H�t�{��@XĜ���T����4�໨(ZTa�|ka�bi���zrϞ=��FA�2����L��L��4�F��1�r,ʯ2�������>��蜝��Mpp��Q\D�'�Y��k�8�M�Aك`�0>��F�egy�=�0A[EWQ�C���Wa��~��c|a�˲'��CO"P��������{��	���(O�C�y���߉���=������P9���M�T?RRA b�3�YA�>BC����T}���0�4gi��LEz�J�|"��LWW��S��UEw��*�o�9�'e޺}�'R������c�B=yx�Sߏg^��
`�s2C�jc�h3�L�+b���Z�L��Κ�!�	��T����������B__������:R��"+�ݷ�1��y:��31� �@l�HM��������w���?7y����4��Nԕ���,�n/�J.))�)ݠ���NI)aӫ���x��v�5���]�e�3�SU,���}h{�����z�y�������1�A�A���} ���WVVFg��1j���X��`?��u$a���:�ہ7cIv�3M.�6H�x��'0�Q|�yF��U�4D�E���`	����i�����<�Gю;����V���(��9�`�P.�����ee��b�-�ey�c�A���8�3
\:66��`�5�G�X��|l���Z�+� Ғ7�iF����������I(�A�>�rNj�@(����u��R�$�]haQ8�k�-~*�0@%�V��vL��h	x�X~���KJ������8^�����Bj�=�[��~k�����^�Co��"_]�@t6����4���՗��)�W�K5���fc�`f�h�Л�ٵ�LR�4�ڛ����3C�w�x�@ر�x�X�L;rV��+� zM�T��'w��˗��9���t�jI9�]z��X#j�(�O��������=L;~r�]�Ә�e��)%��v=�Rx8U�#㸞=��d�@� Rb���^w���%�͏��g3;�p�#c.�-%��(l�Þ<م��+���-��p��O�K�S��$��Đ�Gl���ag'�u �����\O�^D?~�3���C�^��y�������춝��	{�'A��qff�׊���&�ik䋼)qV6��M�������.���`逷�"��\ꄯ��羧!��K3��e g��O{�cW���߬� ua�ʁ�PiA�����v����7X����*:�B��J��yYL3���3��u%Cm���ϥ��W��������:ᗢ~C[�Dr�Ŕ	���iء��,��a�V��z��u���P�s�)�,�P���"�8�.��Ѱlm�0E��c{-����y�g���N�$&��OOK�^{����ma-%�|�ܾ�{��P�M%�`%�2=''��R��E��'���
���F5�Qt�D`���[*r(}G�5�9�%板���,9Q��������P����HQw�4��X��iӢ촐�)�Hd�6��:���D�۠���"[�d�B���`"&M�n���}�������������s]���y�s�s�攚�e �'Nq]�ͳOJJ,�`0V��8�&M��S��wϟyׅA�B���{�H4��}:t2q�5�uu����7﹤�s{��Ś]e�{��~��܋������.�^C�O�ޅ�}���C��?��ߋ�'f��+ݜ�?��
h_�\|��|���,,j�[<�t��F�o��׿���O�P�I�	���
^��OwA�t����"�|V��{xb��i��N��
.�9��]�>~|�}L��-�!g�B�|	����q�����Skk��}�i�������;oL�>D��fU�c���p���"_±g��f��K ֑����޼A���B�I7��ߵy�1���M+�x���s}vh�2��]'!q�̻�|�}JJ�ϟ�rL�o�_
��=��s#Ӳ$��>��$�Dz��mI��p���m�>�:pP��?���.[������~����As�i��+T�Y#`�Ho#�j���/��W�������kfM�Bs4š:7$a�����#ϓΟ���7�Zh�e��?��4Ȩ��>ɱU�
%W�pGY?wh=��WY1̞ff�V\=p:n�=ڱ�н����Id�y��|�zB�L{��$�[/2�t�t��+t�<k��u��eK����A N7{ʰ�) ��`�̥�{+%))��ҩ]]���/aKu��~p���W�*WC��(*)1��={�2-��q��2?��{�n�)�$y�bR��6�h|_�숊>�A,+�mdl�g�Rǩ�b���@��'O>��B���3#�%�����R�"dn���mϐZ$�<L�T���7)�j��><�+�ܵ�ӻH��?ʴ��j��z�/����4$D�	���v�+5ㆇ�;���_U^��ڟ]�A&_��
��gӿC��3����rh
,��>Ϸo�f2�6*NxoLE��Fv�@�8S��,6�[��NU�d�+*5�T�6��Ǿ���쮧�ѩS�������o><��)t/����B�f��-cx��e]OoI9��9��Xwp~��	_M�I�n�);,�<�����3��NΛ(pd���i#�(U5����l/u�cf�)�Axe��Nq�[Y�	���#k(�V�v��\V��ٴ�Pߡi�aYl�b��;3�ЪȕKh��u3�\M��E���χةCZ�_�~���ϒ�`i��/ڢ�t�!eI�?P&���%��̓dOC��n��O�d�]�Ç��� ��T�sI롛7o�}?jQ�~4�<�[�y�҉�CO�6�z�z���Q��FC�����>��=�~�a�;���^g��]�S�~vV�Bt��|�QĆӑ;7[��9�b7�����1�Q�#�I�9g��]��5��ĉ�p����7G�bb�_�Pܱٽ5�3��rc:;{W7c~ݶpv΂B�^ZZ�"��k�Ii�%T?;5�R೑��"�FU���z&;�����bˬb�Yo��>>E69�Vo7���M]BB�_�屚~���y�l(�� sG������%��]���}������\�Bh����EP��rAn�~����""��3-B*m����@dN�U�g��q���P�\h�oim���˽&���T�.�ϖ�H���[�O�Q�ir�h������p�����:��A���R��` 2PRp��682�ao��~����<�ݏ{�5�䷛4��A/�;*�Y���,_��6�/�,dMZt�O�c:����ʭ

L�K�i�:�'���,b����&�S�E>EE�i�Qs�_�L5`�״>2���l���_{��;�TAT��l:u��w���@�uu����N��P����_8|�S�����2�x&���
ܦF�F��]ȍ���H��]_�7�Ե���,R F|懶b��{��rЇ!{��~Gh󈩮����C��_mf���W��|F�<c�~]s����h�p?�W���O��N�������eq���b��5��zǻ��(6����%�$^Y��е�W�F̍Wm^�����q"�H ht���F��X�����U:hB{g<��|{i�z��fDZ�Hy��f��l�r���,���F\O��0vY��/�S3(o�\��\&y�.�Vj��Ϸ��ii���L����/��c��Ɩ��VDPh��
C�Y�l+P��I����ݲf�(��{�U;�<fD����ŴިrZQf�s+t���^=�l�*պ�T|�DMU��Z�,˰n׵�þ}Pୠ��n_=�d�\	}bD�e����I�[x�p�z4[-#--�0S�ٽ�5����3VV�oֻ��m,��,+K�����Wf�9�����g{�f��x� MK���5UUC��^~F�Ӄ�� �4{T��8�� {j���.���_�=���Вl
}u�e�ʯ�,4ڱ�MKK�6��v�J(�˄���p�no�b]ج6����:h55�YU.t��7*kMo��j�x���ܡ(�Lh��jv�N�b�����}zb5�C��>."x]�͒�\�&kkk���y�ed���S0�,g�%�r'ؖ�,��N�N fF���>"~uX�5�kѽf+��Bn�,��5������Jq�,�jr5E:)ŮP9'?���PLD_�Sl�-��J𝬌����nK�,>��ْg?�|��e�������عxv�9�b�%�J�b�@�����0Z�QɅt)-O)�FZ~A�q��MI�������ʗn�]k$����H��;vUGmDS��T��Yi[��"��]�ot�1���Q���*�r�q��Z��\�M=$�g�t[ǌE�agl�����b��������kb�f��+bD�˽���f�ie�EE>+ŇA�Q,U��%[B�|�z��@�������d�-ǾK�p6�[���T��9�|2�on|E�g2)�8�R_���u���!_�[Wӽ�fʍ���WS+$f5���ʻ{� [��	��5��J��+�/;X��~��xz�}�kj*�f�N�H:�;�:�	Z�\�<��=3���/xU�d>�8\O�,�B>э|���0y��jϚe��1���*��N�)0�I t�|%,}��&#s!���T�GQ/�Q����;���\��\,B��ٯ�d8�m6����3�����
~$�W�i���O"	2�c}�g˂��G�$��q����X4�-�l�<�%��|���EƖ�k� 8���_�~��RN����C>m<�B��o����Lb��*9ш�ٝT��	�q�Q���J��ጮ��ж��dߥL%�� ~ii	����\.�=;���?x�(�{�2�������l�x'�`1�Fŗ�f��ƤYE���m����h�tS�K!�tg���#�:��^�,n�����D��v���P�A�
��K=,h�ۀǭ+p�Ӑ�aI��*u�~�q#�G�N�퓏J���jEW;^�M�Hr�K��s{n�J�dv<�R�,:~����s��z��I5���t�.��~��r�
�x0OOŔ�ҋ�L�V�'���dY؟��R�/��������1e���W ?�Ft~5^�����v��Xx3�6�5V 50%��(Χ�꓇$���F5�'��c���%�@�\��G�bl���[�4��8n�9`��jP�El-���p} J����j.�}�����lΪ��S�!�E^2�\Mq�Ʋ0�7+mС����X�%PʺDhU].���ͭ.�gǜ9���-����557w!sg$h����yЕ�뾮9�*fb��.V�&��Kw�6[i���%���Kmħ�B%�vf�3)I�]���~�7��/��+�*/Gr����es���y!��?��;�J�d�y���>ȇ7a��V�BB��+/����S�V�#�}|�fg�9��TYI;i h�D���>,���?n�.yQP ���~aC��_����&�=R��|��*Ò����]J��Gd���L�Vȣ?��.=��}���6��b��w����n���g��تTFC����ujB"K/�i�����G����P{ׯ_?8�hP��^]�^s�Y��?�oH���5�-X�WүX4�h�#���J4�E{����|tl�U5�͐宋Xh��=D��s�F�^rL��l�3 ��PW�+���׋Iayyy�H.�t�X:>P.�Քa6ؠ+�᥼F4L�,�$Z4�Z#�������[�+>{����]�����1j#_XE�)t���G{�#���^���h�2�����^�\
+r�5��?�#:�#4C �h����\yb5�)�zlտ8Ut�T���%��d7Yn4�4�mq��0�볱T	7o��g������3���"��B>�
��j�g�}`;�p'��H�w�����ć��}�QQO� �S�q�p��vW�@˓C��������U>�`^�P�V�!�1�"�*K$ދXB���A|�v�`���^���]Ǭ&q�J��s�����ٹ�����Om9
�.��<�@���=��h ���jAo�[�ԋ����W����ע��T��Ϙ�o�OGhXX�������,'7Wᠹ����\`��3/�1I췟^PRR"��p� �*�F;0vq�7�GD��fc��n�L�`Y����Q� `
�T��>��A#����xQ��DXU�� 
����͍�q@���@p=8��%뢲ɝ��MsS���b9�-AJ"]?kd#>�"����ѝ�j�Z��?ӳހ��YKۅa:`��г"��{����Jk�f�f��q���R���nk��6y,�~��c�xj#Mt`�f�ޏ1<*d���K��C��g�I�h��<�t�P�������U$��ua��0��Te����:��_�ܒ ��ljߜٝX��>V��Z�(Z�X�y�����_�����~vQ�˗������L�JOL��Ҡ�qFd@�C�݆��|�6/o�h�����Mv��l��1�p�
�1�I��6Z�VD�B̵�םxX����DT�f|��I#��r�@�^��y�3r+yK��XA���Nsb&S�2��4,�]A�1B�'�Cۡ�ܮ�213Cڤ�wڋE�pV��ݬ��E���-5�o���9o�9Ya��*��TV�Żv���B���$�pz_��4÷[�+��f���8ͭ�2=�t�����y��g�M���Mn88��.Ls�
�����eB��k����&-���>����,�Zjg��9��!���,��C�`���i����{A���\5%�[�TF`1�CuXk?�/ x]���J���U�9d��f���]=���Í��a���"��-!28��`g�#�0����&g���W��NߛϷ�"�e��&�J���ţMfHJg�N^F>�>b������/���N�!%���uˤ�����[�s�w�::�`���D (!=��v��:&OC��X#�g �E��}}�(�o�'l}D4�j�RW���C�M!��jܐ*��35/��zB�[�T6Q�&����F	T<3����q�=�L��*{�2z!k`�989	ZrB��Sj�c��M��U�[w�M~q�����:��+{R� �Z)c톱�A B�X��Ǥξ��p����xvH��G.��������:}��ę�2��*d�֗�ȤN����W�a�aF}U3pj��_82�Z���-!03��0�e��J�f�;ھ4�I��J&Rg�.N�|�~SI>�	����c���s��A�7�{���ПiQ�Y��0N���|Z1p4�����^�fBZ��6��hbzbx�z[V��܋ə�V�?cR7"���/�rB�taf�ƭUFFF����+C������w58��a!�_��/��N����RȖ�. ӻ���|����A �Ρ����&R�nZ��[�!\�	�eMDx��C������H��E�E1������g�0$�8a�W	��/�]��:�C��k���3NE����xa�Կ�|{W�R�m�߽2,+���(���Č��0:������j��eB�X!� -(_�!��v낏}[����aA:�z.���WW�Rg�R;�H|��ya�o��U���+r�V`o�a��MC���^��V�
YD�b[�ཙ�AY�X�di`Z�͞��������{ȣh���w B�r@�Fŵ1\�O���� G�K$��K|��?��t��X�h����	u(�`�!�Pc�w)Y���s�D�	2���$5��a%>J�VeRHW���G!H�YQo{L�B�R.�g����Ճ���7ЖO��KCw��-�ҡ(��OS��@ 1.ž�R�1&!��)o,�Τ6R��<iYV{	��m�1�@}�H����{��v���T^��:�P�����U�[���@k�Zc��V��<&�_����$7l��p�gU:��a�*�Z��PA���_�DLf��Zo~����{�0� mq5�*[ qM�Kwu��,�������[c��$D�󽁢ET�2-��0&5��}�E�%�l�	�P��b���،��z��h���ҳ϶�C��YM���#B���~uXmd�=�%P�I1,X��|��Xy�"�7�2����BVA#7�i���ۅ�n���?2�
�&6�6I��T���R��s[�?�
���T���Ŵow���J�����Y8v��p!�֗�{:�Y~&��5�6��06�V��}�-��+�I���Q�������s��;N\zCsy��d���߭=�oρ�����!�ϙ���QV'���6{&��c���㥁 ��݉��"U��\j����ˣ�!&n�`��oe�@˽?N�a�I�/QD'�@A�s/�Eh0O��{8,�t�������T
����j/4xX�i0�=�)��;��mr>LZ@xK�ݡ�`5ǃ�B��<U� g�󓰻�84� W�B֝���s�%O��s��w"��{��r���!���>�i{y��V�!��W�F��a�L>�>MK&^؈n���zM��~T�ݣ� �Zh�a�9��=�T�]$<#��\�{�RJE�����!��P>����U�9��$.�F����c�md�Tll=�AQ���zx1�a*��'�>�<#U�<�����r��{�zH�J��>B�~�p�/�"���r���������@��w�W��pؗ���o}Rԃ}�6���8��IdxσyZ��|�����_�kYs}O��Q߁�ۭ���)�~3��H�/XB�v�.V���{>{o#��#%z�סd�`������6����?3��BJJ4\��O줔#�X�I�=�@	�6A���Y(�����7��ӚJZR%�)iis��^�!����S�*PwU6���x>�})V����|1��rix�9���z��(J����-�0W��b!c�R��J3<����3 psMo�#4�t �۞d��m�Sf!��XAyP�����<G=�B|!���E��_Le�6�=Fhm��������e��E����=��{y��c��������Qb�o��掦�cr8��|��Gx	٫j�2������V�Q8��rU��w�W�(-�/���E���=�@0��^AE�@��(�e�0����¨	0;�7o��0<\�� U0��\��5�!(���N���-�����PT�E�=�B|�*�Y��Y_�������h_�J�Gf2m���u�x'8 �l&.�
�V.�ɧ���\�)^ (-�ּ�������F���^Ed����O}��V3*:����w�"��l������\uW]U �	/,1� �S�Q]��b	x��M���R>h���9�KvWk��U@c����ۄ�y���Mqɓ���ˈ~L^TT4ΑO��[���-�ar���PQ�	@dlT�@�KE���fm�3|	i������x���T���;)�V�@�WP �a�H��!j�P����"���e9�Y��ɿ�e��JONK�G��j�Q��3[Ξ����z���� ��/Bh�&�"'�*6�e_[Ȣޅbƀf�r��O4{ ����ٖ�j�s�Wj�mZ`$a�G������$��p��#ڮ5��oϤ���$���&�s1m
�q�]�O�.��� ��ٳʿ��\��g�� ǯ���^���\�9P��X4�,�$��[N��E3 ���V��!\�Ҷ��*&uˢ�?w�4�A��,ּ����ݖO}�1ߑ��+,؀�|��͚����u��r`T����OV
.  ���Ѫ�u���\��o���|���^�#"U5ፗz8�H�(��g����,��^A,1jF���DZ<�<�0J�1	�7M\0���<V��ym{נ2ς�b��FF:sA��,)���,?��� �N��OӶB';�T[C�y,0�}[�&'���<��d�XHY��,��ZB�*(���+�7b6� u[��%r�6����~+wQ�d��f�ӷ��ʃ8,� �j�;78O'fK��, X�L�����C���?�E�nw~�"��#B}&�&?�0]C��d���']�q�1����V �^{Zw��Ql����z�w��B:��(
,������!����'�Bl�
��e1�<���,�£���ַp �``�^�푆%�=,t-��nf~��R���"�K��9`�[��%4�v"����D�	i��ُ m�K�����N��~!PP52�F�v���r�5�FǢ���E�
O�H�pl b��F����5�@�f!x 	�Y ���fH����	��* G@S�b�-(v�ᒁ{R�?5%DDm؈����A���&3��[P��%@�Q�I�%�� �,�.Q(_��w *	c��EA)�k�>��S]��⊢?E���o=���2U�nOJ�+��z{H'=m
Lbʍ�E�؞�y���7S�P�A�n׉��k�\�-!���P%�D���S�� &�"&���_'}<��]1�$}�*�Aޖ�pi%�t$�$�b���>�,d�qEO$7H_U; '�ٽ�{]��5�7��+܀~�O½p�Y�W�p�/�#,m��Y++_�'4s�@����s��Cք��!F��KKS��޵F��S:�
������G�7��"�S���eEb��PD�Vpm�Ij��,�Zw�.��u?E�,�/E�d2g����L��-7�n���P�b'b�)�"pX��"�け�Ra[�̶�Gܼ��{۞� ��'��hP�ٓ|Gί��c�Sߦ�w!�n���5�/��f:�4�V/��#�٫!��]�?ձZ�['���� <��+�*K�K4��BJ�QQtfvfi��~Q�?���n�1�̜y��F�޸�&0~j���5%�.tp��`N:\Pvl��%��Np�U�r�".���%�R�1����Z�U,a��7m�_�����L��ۨ��̊>F��h�hK�OS@�UH�N��N�8��Gf5Qг�tY�&�I(ݳ��xm@����������Npf����t�6o(ż�PX̿)�Ǣ�|/A�@�����B��hy�'�7���_L���"�� ��D<�w���͎�>�`n�%�Z���p��}����uut,Ü<|�Ù�!zT6Z��Ӛ�XD��"F��Q�FA����B�=p�^��=�@�NN�ߗL����:��m��<��psԹ��;�v����0���;[�k��;��)of��H
oN���1@��3�<+����<�n�o �<��3�tͳ+n�����)����4������?h�ߔ�M��Ԕ���vi��49�����bn��N������:�<������m7%Ο������o��/M)�·��*50��p0�^c��^>
W}��{�C�����Х�.d�����"99٫jO)'xw{~����}������1��C?�#�,^~�<����	~�GUph��ck���ח.]o�̓�:5�}!��G��%���em�GS�SN���ܜ0V��Y��gZ(��gu$�T4�M��%>���]��9.��GA�}�h���v坾��YB{�v��W�B��c�������~cᨁrҡ�16�-���'�,��1��6MZ��{<������ڼ�Q�?���>ބ��?�3(�稷��N���x#������`�k�k�����8H���U393k��D�XL{���;t!�2��6��x�3��G�Y�͛����Д�n��w�4��O�%n3��J��|*�u��v�C��L�4y�}R�w�(�K���\��-�wԋ�&��tV6������Ŵ�OI2|1yO$A�|S}��7a1�x�W��,���Q�&�חx>#�
[�O�7a����.��df�I	�����͙S.ڟ��2��{2��X�ЩX?/���Us�J��bӝx"��?_�7����� O:�t�k�E�����|�}�R�D�~
�S���?
���(XL֋vށ]��~��%�����ze��N���3�C˿<DN�^~n�m"�u�o���2���ny������kGd��y��Ky7��?�J�����?���g��_<=�kk��ԄD8� �>�SQ�	?��E��uM#�\��}�� J������)����wZ�o��ۏK
��x����8r��Lv9#�+_��ZB�]��PP�m�ޡ���D�c`�������Ңh�)w�ܒZиvA�a�$�?�%���.d�W&����ʫj	�bX�y���ff�@�V#�$�X�eBƲ���Ft�T��1���NyJ�*%�N�>I����E0�^,&�}��?z�iwKEpt��� �q�l�3?<<�vtr*��= 0^�q	B��u����o�����.���r>����q7���,������7u,ڌO5������Q��c��/�P[�A���Q�d��HUB�?���t���*A������L]~;��wh�h���x\��ܼ}֔V�8��t'�Wj_XU�$!K�e����%/3V �˯;&��A�ǧ�6a1
y|�v���ڻy�~����n��sU�b��_�M/�iiq��"}��7˿ՠ]��[�8�ay�̕�Q�1�/�H�t>���!�Qj�Ӛ���}@���os�ip����2�Y��������F��>�n�Y(�Ï�Vp^���`@`FYoT"W-衆�`�����i{���x��r4-��9ދ]�rO�l�-���s&�����du]zެ?���z1���a꧂�"��I���~�d��2^RT]�n6s���zM-Ai]��#5|lGq�����r�^� N�(���#��ި�H0˝={���wI{Dy�d���Ӽ��#ɶ��%��^-a���l�J� ������8,�J�Em�6�n�DM�4�t̜�n��>�P��:�5m�����D�KА!�B����u�)�}-���T~=~��U�ߠ$���_L!��S�5i�%P0*t��G��D*e%:��E㪷���_�y�߾ ��BZS��&�/������tQh	�J^SVYЉ�k
���x5���ua������'�wp�1� �Ŵ�Gɤ�����.gXٗ��!:w�Y�[q�xϾ�W"���K�a`�u`��`�,�
%~��ؔ�6��_��+��_�~�~n���]�z�,//�9gi�hևf���,ֿ;.F�[sY��{z���B�I;SS�� {{�g��%�Ѵȥ눃�c^��q����o!^8...��˯�B�β�����;��F3_[��zG��Ƿ�]�G�ߓ#x����g�PЫ�0��#2zz���A�6�� �\���55���f.[�
zC���Z�#��`p'��9��a�1y���I��yMj�J�i_���N�[�p�g�g�-d�Z'jiWD��Y���Lr�r�z�Z}Uͧ�4��o���΋Q�/zc�'&&:B���a�����(-�}ݛi�ҕL���V8���3��i݂��v=ƀ��n7Xv$K��̉ϱ�U0V�ēL��V�EeƟ#�SA�Nv��֨&��5������N�|��/5�i�kwuԶ���ZV_��6Ô5x/|!b�;�F|�A��^Y���S4%��gS�A~0ӺX�4���=p�pi�=���0�����e&� �TO���t !�Y��t��i��$�LVv�qb��G��G�î�=�C� �>�lr��������|�4�F[�,���5w��yjTXT�vw�yvW�R�R��6����e�wvc@����NiM�`ɐ7q��IȆƞ��23�h���ր�f�����gr-�g�AU�9�aG�c ���+���v@��h1�ѝ��3��U=��H�S���!C�X*�9���/�Lc�@Y�&�X�W���U���I�}��ZZZB�
_s/vuV�f0P(�섩AV}z�y~y| Xk��7�͵Y�CXd�*䁣�YH���=}�`�55�J�@���ҫS�~S��I���U��č�y�<i��1�i^�;�g�5�5T�83.f��6М8����hݳݛ��5X)�<����L�t��q>}8,Z��5�kbi�^�CM@�ib��K�&�cl�܆��0d"M���f��ԅ�����V����V�2�u��+a鹝Ú�D��� �	����>9�o^���5X��������N�5���D��ּ;���6�*ÜU��0%��u��.�hfV^��?�)Us�ҥK�>-P����|+QQ*n��7c	�u4D���0��Q��Ty��h��Ma���j�_y���Ȟ�9�����?�%��X��%�ld
u��>����ߍ"�~�7�!Xs��8U�']�>�>��q3N�=3Ů�ג՚�'�P=wl�^�����xX߼�{T�߀.B}�$/slj�,�4y/=�L���E]K+`�L�e@NϚ��Ԯܤ�g�2G��t!�D>�^6p5^�_���~�2:�3Ͱur�]i�JN��N!�>�<�L���oAB�����&Cw��Q�2tْ�SX8������L���ʛ�6,�'6�]��q�t;�^7X%p��u6ͭ���HSd��/��b��q�:gz9Z,�[��l��w��MK�6�H-!�H��1:��؆��I+WK����)-���z)/l-T��f�l^�vIc���� �,�
�;у�� �&{�)N���5Qtu#�¢����X2�N}�gw!{H*++�}�}�A�@V�'C�<`<����3�JʾX�b����2=>��
_��d��B��>}���S��ѬQ��Ǥ!{�K���N��k��֣< �=��ƐH#G����).�ye�I�[����KQ�~�6q��S̵TI�M�	�����~	`� ��C��_Z��<{���Y �];�^mМ�(�JK}����`�X�E�p����m<w`h�U}�G�܁��Ԥ�;����-=== `�$��6��s�������s��}@�3=n�'�~���uX*`z�{
���2Q �^G����(���$,�F6B�#Ѐ����.C��5�EY��M����&|�U�I��)h𩏣pӄ�]��W�����Eݟ��W8����?�O��F4���A��(Ih������(7�.�2��P#���PY����2�׳�>l��W��!�F�ͽ�(��3�	��k��¦E]�_�~��u���+}��1\l�t^m��ҷ�(�䬲�1V�>�ϵ���n?{z��C��p�V�����7�Q�r+0��r��3����a&�9�rZ�OB;�c_c��H��-%y�w��߷�~Oc��AF
E�P�`=L�ꃶ��"�څ�N�0�Y��{���[��������m����n/ŷ:�ܱb����ML~%�pp������(��[�˺��Rʍ^8�Xi��Q�5��C��%�%^C�I�j(�@�J�12�������(�}���!��-k�K���mɟ��-��W�@�I�hF4hf���
�.�TT�C=��$��Q�ԀV�k��F�R� �}S�
� ���m1�f���V�t_�$
/A��Ð��9�L�)��n���[��IHJ~�G�]�g�ÈW��S�)���^{�OЃ���P����")3c�`A�tK[��T��/L�ϩ��p�rBMM-OE�P��1�҂�YF�6m�<3��z`}�rXߚe4�rQ�V}9��9�s
_uv/��j���Hp��ڂ����gA��c�jΙ"�2Q��UfM�����AG��e;x�(Q�~��*�6AD�Km"�']�̍���6fU��P݄�1�sz�d��k�5��@���j��=�U�dV�摻vU%@EWCĈLi��h�?�	7����2��
�V��1=�Ll�ѯ��V�ڲg��j��TR2�c�4Zw�<^�PqK�ak��O��>��ҟ�ּ�
����u�����e
2�'�l�$�4�?�9Y$ؔ ��VVF�8�Y��o�}�Xt��l2B��Tq|*�G�/Ͼ����K��5ss����.�ӌC�D���@��t�*[	��hǾ�|g��!�$�O^������I��W �,�$U�$��/����r��O�}��f�|v�g����Q�@�(�G��u�-Wj�������}��h�k�Ǧ\��{�� UN@�;�tkS����^U�L���O����
�f�ZWf^$�?
ι�b�
'N�;��'�Al���.�q:=F���߃fc9�KTϹ0\��t�ji���|�@�q�ӂ���;��s��� A��ck)��a~'Tɓ�پ�>}"_�@��bS&������1lT��W���XL�:�$���e�X��d�j)L�ٱ��}ך��2�!ٹ�1cu+��'i<����<�T��~�����i��lG� i�ް(���/���`���R&r��08g$*Ůt�L��w���� � ^�p�e��c,8?c�ax>�Pk�|%�*�&7��؜Q[��9�'�>���v�'�]��sI�Af�[���Db;��B>�px�I
I�k��q 7NE���%}�˯@�(\a�c+��Sؚ.R�A��}�"�/
��'���}�h!�Ѷs{�\ў�����2��ln�Z`=����h��
tғ6�Zq�$W�%��h���7����Ӛ/��)�%��צ����dZ�~{}c8�p`�K�]l�L�+�����"��~=��u� ��i��t���â�r�p�l�j��t��V$��R�~<�*�Ni�����® fMߋ�����׭���K��T+���O��Zd'c��-�	�����n��3��JNf}��kOk����m�n��-hj��hv�JY1iȍ���� ����S��5���{/�9�N�
�D-Qa��T<�\��ZF;&!!q<����-"��Ϛ�XL�cz:�A����B*Z�ZC[������{���l��#dZu8�0�D$�m=��e����k#�T��M"R�p�!R
p�z@<+>�xӍ��I⿽�h�H�H�f,ӹ^���S�h&@3�N� ��k��ӕ�'�[�9�	����@]���S�<p��x��^�1�/��/��K
�ӽ��'�)K	��7Z^�ӻ?�Oo��P\ʕ��n�̶�ї�Fo���+��O�Q�,sb��<]d}4c���A�p"ǄO�p3Lw�k]��LO�Y ���ȩnu
Db�S�!�~$�;NUM������n�Ѥ��/�b3@�<~���mڨ�6_E v�H���N�2�^�k�؇�?� r�6�F_g��ޝ|d!�:�5��bGbG�?lA4F���1�����u��4o8-��
���L���	��EsI�c�t����`�=z�ś������ϻA&���L���-���l�!���Lgf�^��ͼG=�e���I9U2��M����:�,(�|Q���.�[�a�ID�'͎��r�$�W�/]���]��j��fS�u�E���P%Mz�9�������l�N�.�Y8�q�\��U5�����0�s��&��_�?�N��^��&� 0��IS�|�6�7{��]��Z�d�N��k?55UJLz�j�Q�3~���1,#���E|�i!�H۠³y�ORAȞ�V̳�߃�LQ���U'ARކڦ�����p��kEH�@�m����+�zj���ܾ7�(�G�+8�C����ҪFE��>ݛt1ݣ*��� �Q��'��i���deHr��@V-�ܱ��z�Z��2�ո����Ya��E����Wt�P2�Rj����.��|���h��eT��r�&c����X����i.""�%^��ޝ�ƛ�H�A{~�6�3�g
�z����A�G�m�9<'����h�����-��YK,p��P7!��� S��{� >$�[�=c�㉤�bQ�o���+�x��TV�`��d�����	��(�u���vq&���2�+��Ϻ�h&⪨�ʞ������
�tO7j�xq��>�쏄8����u�k���~nE̋�y������ q�������J�DYFW��f7���~��s躛ڳ/��S7�J ��F�z,�B��Y�R����B��"?��\�j#���{=h�ǻ�i���d�Z�Md��IY���f��=�e[eJ���O$�h�Z�����3������g��?�=��d򀊺�ff���K<f�*p�юաVέc�ЃZ��|�;��a����4���ܢ���20�̜�~vY������N���!7�<�Q7�8��};"qޞ��>>����t3pX�8�R{��4OQj7L��xT3z�_�8�g���s u�h;Cy
�[�m7^�{cl|��#����}x��S��VE��.��<���B.�}��Jl֩Hs�\��Ɋ *Ԩh��BeB\�,UaD0���-��DkY�B�����s�{��T`i�v�?n�D>"z�	�8A&}\
��Rl�1�B�.H��� ǘ�6n3zp�/u�E�X
�bE�4��>��~�J�
cX�1�䞟���b��:�',@��s�z��1}WMЭе�9*>�)�=7�	t�3Ʌx	0���K�c�*Z;�#���}�
؎}�2�VW&Ϙ.ӭ8۷!��]��Q9�B�T*+N	����qjp���83W��ّ ~ϓC�/�Kr.�7��!�O�w�R�d�dq����}����&ɥrxɲ�h�УQܕVH}E���T�eLגIj2�zP��������v��l���
CI��"|,L�M����Lf�%p���6�Dg �w��5��0kɟ� �.C��@� A��
��)qk֥��"�$����jg�@��#y��I:4���Y�Ā� *2�ھ�^��� _\H��� ���j��U5���
#�61����� ��M&iI�2$�w`���V�I-�J�� �LR�����%$�Q�I��޵�`����<���NB���ND�0Z���ǭ�	d��n@�֏��I�k�͞�t�kW�g���Xu��_����j0�b��:�F�����K�4�#���T���mܯ�<x����#���2�`Ц����?Ae]@�����\�}�o�S���!G����
� r�����]܂Ԩ;T	,��6m�B^spO	ZY�m�n�, }�f�}	�{�H�w����ߖ������!����D��f/i�Z��b���f��(��ϗG�H����VAB��ln���%�?���뵸����@�b���9ovJ�N��䑞n�	���Ϋ��T�$}���� �W���܋e٤!�XI�B�H���S��ЃM�q%9inE&_��\��uF|�^�?�����i�'_�nuvH�+Ю0��X�.TA�B'� Ө5��H�"�VTTd�^$x��vŰl�;#�S��I����Cq]��jB�U��k�q��f�! ��t��wO��T����a2��Sa�v�k95]�`&�5�Ї1<�p�⹫���+���]�&�G�����B����{x�k�L���c�-�.*����[�X�RzC�����V�Nh���yQVƁ a
��b��ќ�b(�IG�pX��;�b������e�q�"٥�1mRh�ź�����,���eJ��h���%
���}�,���vq.�����q��wR�B�J�h4�	�}Z�WO[��)�Ľ[�� r��T�`1�8
��[��P�!�ֳ:�N}q.��J�OԘ"���C�:��H&E�}dlL6�y�E���������/pj�L{��s]T�m@O��rE�+�e:�bf��!���<��4�8oSm_;m�2Л�Ye�'�L�-�}'`{c��S�wyYp#��*j�*&�j�/�!��9WLw�l�S�� �1,� ��
3��j�$�Ǿ�c�SQ��-@��i�n"��%�_j�(3�N����xiKX�J;���`L��!hOv2������m333
��Ѹ�� ��8o,��]�Ӎ��]0�ڿt+�]�&����|��zt+z�74����J���h�G��� }L=�I�I��޵&�l�9i+Y]1�^:d�RTxhX�� ��lgr�t�z�Q��� y�����T��c�Z`���d�"�b�C�E���u��
�'*���N�TD�Oa�Q��!�t��?�S?͢t���u��g�Z$�E��f�'�橡�G ��w�X*�,'_�����a��u�p���B�2����-�O$rI��s��(j��DL����J���9�CN�E=����)���{,�`���B��
���g=;���w���K_?A��3��t����d�弐L�~7[b����畗CH�N�¥J5�ȋ&U�&�\\�&L�Pe���҈$X����4����?D�vi��U�4���!�APA�%a��
���	�q��+�"� Р� � F�$�������eWM�TMM��?4���}��s�Kr�<��ƠM��'2���=W��!������ku�X;u9ߠ �o�5:i����Ѭܢ"�)cSj�9p\#�z��o9�e��,�ވ::4T�*�$�'�������_�LhV�+��97>42�f)	uq�����`������2hP
AE������ӵX�9�\�`�ms�O'�To����.��K`�.֭�ov�B�5z���:47�����m��|�CRe�"-�G�4=8%L|h� )*�D�ۡ�r�Rhe-�"��"݁�	�333�����_���^�Ű6+�F� X�"���O���D�Ͼ��~i09`M�c��c���n)���4p���6i�u���KR���T��y^3u�AcڍB܅��s������C��{?}RO��O�s�h���P�e�W�As;'�U��T�n��Ƴ��<H'�it�t�;���X�;��t����Gտ���S���-Po:�w��\����I�o@3�9�ϟ�=�j�-�8+�)ڦyS�]�-��|dg�
v~1��|i`F�mJ��Fe)g��}� �4�~���L�X��5��x��-����XJ`���d�jO���b���&-D3P��I"~L��g4�vd]��o�(��Y�� nL~��'H*�;�������|��ZO����SÐ��*�E��u ���~�߇�
� �J(f���޵1I#���i��4w	�[7�:�ʬ��r��Խf2�q�!z|p��+"�Aޡ��'��Z]]��5���I��^}ceip(�����6r$�W�Y��C���i98=����i��~��Pcj���	��"�����b]��&�q+��b�G�;I�`�H��9֎�*��Z�E�����!�<�B]_�W��S�066vy~��i�_�6V�?�fИ�Zo��gǳa����(~� �RHP�����t*�\��$�t5��ѸKpX0�)�?��]֜[	�3L����7��|9�µ���_052�5���B&h�'�M��}η�N�b�Wśf�1j�f �C���Q),�DK��@	��g���^���M���*Ć;)p���v�u���P�,�\�s��^@��|�������k����###��'4F���G����~�Ih���b�ξ��2���n86��k]�(����=�N��m�7XgD�2{�^�*��-��<�}�W?��UaO�}���4T����ƿ�`X� ���l����KGڵ���&>��X�`;;a��\qE]�_oc/�A*�ŀ[	G����9(]#��w�V2p'�qP�;�h_�]�n�>\)<\W1[%�yҮ�hX���^#��Δ���A�{�;��p�v�-���֚h:��.����!�;0�*뤣����S�r������j&���V�w�^�	܊�U���\��@�o����܄,� �9�/5U��uu��v&��ָY\�t����W�#�l�a��gw��ЖR޳� ��+���l�h,|�7<	�Z�x�~~��O���G �k�~ɣ��AX/FjdEc�;�[>K������[���4+HC@�P)��Z���!��Y���*;�	�tPRw���[�|�����m��v�1>�F"5��0C�_g��2S���-��rK�☽ٔ�rIP��ל���9M�R p�@�n�ؿW�f��{�bF���Z���~:8���xI^����[�M w����!�W'�!���O琤��Ҽ-�s�3��S��|�.���
��g�NR�|;8�� ZOD��.��[�Ei��P:�k��=&,EͿ����5��(T����`����T�POiI�ͥ:��L#���� D`�V�&�+qde��U�1t52*w���� �E/�(�DO>�m�U� ��nS�°���R�6I�nC(��w��e��ޭ��3K�`�b���������}�0l��_��������t�jw�?�!���}C~���t�Ƙb��K���4�Ǻ���/:�3���vCq��'�.��7��p���m��+W59-�>0��æ�ˉ�r^�ƫ��䃶����I�P�����0�Έg���������f��?��{��j:z�o�[�.�V�#���aNat�4V����J��4�n��c�rg�Vl�� ?%�[�=(^�IƜ4� Wq������I,����[ 
���y� a�I��	���b�z׭f���+�CK�C���y���X��@�DvV���d�q�~{�4B#]"yټ�d���6�5\~3^�Ix�Y"2��i�0��GK6S�l�n4��:�E��L@P��d֬_�҃A3>j(�����1�}��İ�� �, �Z�~X��w'���hc4���(�{���_�U����\3���n�+aN�p�.��f��N�L���!g���.��3�\�5U��A�����deА��T.��~���D���͌���^,�����XY��f�����%�/R (*j��FW�Fs���`�=������l����3(#%`(tC�G)��\��lx"v?N_�V�9GP�X){rk�dq^fT��d���X>�c ��'X�0�Þ����fH5��e�3�H_��cT���R��ߓÌx�:��8����V#�����Eu��~��,��`��@0���n��[�^���m&�*l��~y֪�pp�������L<~��_�P?
xw��*�@nb�� 5-+��	x�\wO�+��g,�Rb���	
**���C�~���(�2����5��"c;��*����	C�#������`��P�	)_�Ic-��b�?���ک�j�ik� ;k�6�@kn4����Ϗa�,1�cb�1,���c��MZs�ʧU�ޜP4!^���w�Lԥ���q�}�ꕒ�/�[��0gDA!�p"{E�?��N�s2)�Q#��ɾ�}[��s[��ꩆ��id2�5QZ��,�,�����N�Th	�p����T�$`�Z��fs�e�P.�4�ɫ~���@/��nU����ۉL�E�se�F���7I��`,_���z��Uׂ�Rv�ZYQs���=�K�˄V�~�L�;��̊�����'CmY�"_C��w̆˷��	'�Qo���F���_����+,*��Q5�X5���Fw8�J�''&�� .켷�(�Q�	�,����9Ws;.W���1��K�9&5E�,�ј��}��{�wY���&~+���G�H!͹��>ju��+n�a4_�̄w�����s&�&��'��u�x�~���-���@0�[����Ɗ�5P:bJ�LfJD���d�n���T���N\r6�?z5fԾ����רg����W�P�0�/Ϙ"�u����x��v�M��Z$H���lBxtw�J�r���K�M��1��<�1�U855�B5�Ue�Q'�7��{c�~@�6��@f_M��;��nM�&i�[)JW~�2(��z�oO�����rB������ܢ�mB<�hѷs�o�?D�!�����DϪ3��Y
{Ҝ���������	��_C��۵(�[��$0�?	^��R�T�uj��>�M�?Do֭�oÍW���%;�?B�wxdY�lo�|qT3���5��]<�R�~��sq��,
��o]]��5H�W�'=��3�3�ڄ4h��.����TtQsmaw�N�/[�s�+�L콣���� E��R&g���I�?�NI�_m��OK�:Ύ����D�+�$�lHY�<<�菮�e '^�NO1��/V�0O"����yၫ {��٤R�د����<�K���~�t�A�W-�i�i�-e�F�t��ϑa+�Y��X�	H8ƟW���݇�B��ZG +�Y�8� 8ߪE�{�xn]�[+�����c!����ƙj+Ʊ½v��0F2j��9��q�y�F���ɣ8F��#&�[�)l)��\F'`�j�-==}�+���yCaa!g�]�l�3�\~�����#V��W��EEE���.�m�x�R���&�U���;�/�p(%7�%���ӺaY��RGH��K��m��K�4�芨M����O#�uz1�c��;3Ir�n�R�L5��rnr6,zwZ�����ɧ�s���ׄ��F,���mhh�aMԝ�-���fo4˲��U�{K�+,���[�B�fgg3�j�Ǚ��m�/��	�\�<<b;v��N�g��'�+%��"q+:�ӹ���L�Է���s�g;!j�]�s�C��������58Ty��}�_�j�Фo.��w�k%w�41�iM�V�n����զe]Fg��������#=!��"�]ᠡ��X�Z��/�.ۮ���m$��c������(Z
5_�Z��wu�}��ZQ�C��{�N�����r2�����P��fF~p(AES�'Jς`^���i!ƃ��?�%$r���+�R�� $%�����h��5���Ԭ+���P�w��=���C��t.���ּ�&6N�vUD�c>J0wʂ�M�Wg6}j,�f�|6�u
�͞:���"Ӱ�<�-�Nɯ;��N�%P<P��.�B��Z�-��Ѭ D�o����	��y��6��4�D��a�iC	�Ncp۝����J��8Дc��6���eV0D��؃�y�s�?�{����V|�h3�-���t�v���$��Ӝ���6��ey�����%���^�v�q��V��S޼y�֢ڰ��3o�i 
�@M��|�-�P���t*�����)����a\(:����NBb�H�)��w"DQ���s��jP��rwK��������%>�r��L��z0�F��6�y�|�Gz#�%hf�0�Y�FJ9�y��Ǖ�����z�ޮ�%<z�8��4��)��:�����-�Se(�w��r�ՓO]�D%�,�����mp�p�U{#�EE��Y'�}����3X�x�C-?�4M�s���᎗q�X�?*ydEZ�f���_, $��������E�*;׳�7��7�y���~~_�F����Sc����T�N ��� ����Ӿ>`�X���'������J��TU����&�������k���(����}�&9{�.�'PK   �}rZ��g  n  /   images/f636b928-3cee-4f31-b55b-93d56e3d5b88.png�xUP�u��{�;�)�AZ����C�I)�-����8��P��+�{���tw��Μ93�pfv�,B��*�  ԠJ��&��q��un���j�	 0�����z�Hj/�w^z��^�V6 ___>GOk+7>W��S) ��AMI^�/�$���Ġu����������1�6�b���w ����(:��9�A�B`hz/�抉���T�K����%U�0�2!54����+|������#�lI�)���ŶE��V�c����m+�h�@.�����9UF�*o�@��Qt&��t�t�DA:2�L��K�H�e0�j8"0��h�����A�a��/�b�V�D�o��휞�H���l	}� }L�~���>��t����|f?�Y�����0)�){��`��o5����1�䩩��-��&�{�6�P��54v�J*c�?Ν/�yޣ���;_�����WF��� �z����ܻ���1)�?�n��9[��j��U�Ҫ|[;9�K:�D"�m�R����7 쟟[�ެ�68��<Sic�"�lM��ljn6b:m�&L��}�pj�������\����ֶJ�U5�tޢL���n�l�)�ox;nx�TY �J��y�I�@��y?E�ʯ���zZ�Ҍ�w�;��T)�?'Q�63�������W��:�@��e���4�R�I`��V��ʿ׋[��^��FS��'kc��������k����$C��7HY�T���H�"n���v+k)6���2�& �gg���;�>=�y������SAJP��f,����ׯZ�:஀[�?�q���Ǚ�UGtY
~s��^�F)O�\��Ý.�`{��3��b�$�[��H�:/7(���D��Y4�zV����;�r�w�Jtw��t��iYuI��>~ɺ��%�^4%����o}�͊��!b���k����PP�N�˺���y^�i���	?	�<��횇
���<疗9ϺN�s���Y�S�nF��r4J[���松>���]!faU����3�:ːG�q_�
���?�君���g��fٮ��v*�	���P�������)��Wic1�&��
�*�QB�#}�,���Jt��Ut6�c�Y�RY����m7�dgF����w�9f`z~���������4�)�n2~��m������遡`W���g'�x���!���+�y��Dx���/ǚ솎q��0�ط��S�<�+�/@� J��,jnn6�FB�YW�1�z���0i��,[����zUiQ;�D���ϽL���HN[��|o�����\m���UU����@�Q�������g�3Y@�/���Xޏ�w;�s�n�%߷�WtMfI�0�c�IUr�{��K�����a�u:S�a�n|�IY��ARĈՈ�:� ����;4�JMP�64���g �6\]a~��u��E��5M�e)����N;�Y���@̬�{V��ɫd}<,�� rp��!wL]ה��V��`�|��L&�E��LJSKy� ��V�;/�w#����(�.��o�L*��P�,���L��f���n*��/f����k�M��C�I��V�{��f�9��e��x�Wڜ{A���S�z�}������:L��3�DR���5s���l��x9�o!�b��9�!��9�����ӖJ#v�2w48SݷwӤ�Y��VL�kR��NX�I��w�L��/�����}��ͧ���^��hx��x��|Ԗ�+�鳵�	��H|:Cu��*Z��j?|8c�{�|N�1)���.LCCSu����L���(���(]�:��@-�/!�7�?�X��M�-�p�.Jjߺ$�s/ls͂��Eg��L�8�:�?���{t	)�|��V�~ܟ�����n��Lu	�gAOB�����Դ��>
�g���xԂ屙�WȖ ��#�!��{�8ğ]�7�F�G}^���8�xڎV+/��f�}�X��}�,�<cj{h,j���~f��gi��Z�陟�`�c@�3��8���`̂܇�7�7+R)wQ6����"z���:�*��F��7�|l���nI�o;u	%�_�ۛ�?>܃�Ѩ&~�	 ��:#K��6
n�F���4epftg��(���Қe��M�o�#�a��%�:$�O(���SH\'dn��DN�O�)�Y��"<����?c�Ǫ���	Y��;���ª;�lH(�)x[t"�"G��<��㬖�r®�k0�&�`��C.�"0��<e���a��@�^�c��",N<�s�9q x���f�\WOL�F����j�&l�f� �����0����=�����	�@L�6Y�Ed��Cy]���N��5?'?_���Y�q|N!u�ʜ�s��u�N`}���$~��g��^�z�qr	J^b�e�T���ouVT6 R �zynZ�e���ۅ(�0���ȗ�<Y�/�hm�K6`ϓ'�L4a4��{�щO����������"�M��8�;>������m+2/�O������2xS_:x���S���P��A$�޳�l�ϞY�(���5��l���M�'ק*������w�}�����Zq(㪯��ϣ�,�݄1��-����E�w�>�k�O��$ܗC�@x�j�]��O��'N�TY���"\���Q��K�iJ�y��1��欎|��q��b�ӽ�#W��T�Q��ݪ�6�E�#g}v�\|)&�Π��!��S�y���k��i�$��f�*����˫"T]P2 Ȧ��$-t8�j�QG �7��XV��#�{��L�v�&g|�|�;I�Q+>T�f�b�+��s.�	�]t�ۃ�cm]N�û8��z���׈0=XX���8l����=�]��x9��^$9�m��r��/���Ɗ(Nwn��X���Ea��z/�ejǫy&�G�A�1��u^�U���e�Rv��	A���L$��t���k󴊧b`�x�`�`m�c�[m|�q����%�`���tl&i��{CwC�W���v��3zB��/�0
�}���j�FχY�e��QeUNh/�e�违:����y��',�[`�Є���l�#�w�-ܳ�ע�yRx�DE�����.B��l<զ�	�b(Ι�O���5i�K��Վ���R�'C�2��Ut��v���R-�U���H��Sh��W�\h�a3Kf"!N�PyMlOB��	��ɦ��T~��p����&��.��`�|S�����YP�H9B��7���'67���!�2RT��l�K>P�����F۞)/���� y�I���I� ݺ�
혷7������v���4��YH��V~8�(�y�E�l#� ߄ϲ�̲�'7@�eV�M �:P�����D���U9&��*(h���p��`�V������Z��ڎ@����Wu���T�xhT� � �ɣ����w|��n�X����7��`���PI�l�� ���}�wd��.�Dj�z�P�1�sB���E�!w���Q�(�����z�Y���H��-S+����D�Gb1N;h	���4A���	��73o��Z/	[)*�PV�"6ӱ1S�$RϠV�+��_��A�>��2;DU�l��
r'F����m��;d�7V�+�YW�H����4��5K�/���z:©��/ؐ�O��n�w���f�eD��<}�?�Ҽ��_)��dz����"��Y(v�+cZ%,�`�UH��(4���ٯ�P�e�+�靑A*&�4Xf�%�#��#�(�C Tq�j�YSu*r.������K�<>5W179>G��gf^~�Xݹ��������.+Ը�.��� �	Y&Ic0mu�]��;LlV���ֆ]2a.�|�K�FE[o=�a4�X85�=�%�P����V/AK�Ndb$���
���(2�R��t�b������ޜ��R�~�kbs�ۦ�]�{��&S��Rk\B\c��#��o��x��cK�\ۖ�1̥܊ou��p�rZȠ�xu	焝��9ȟާ�F��|nG|Wo�bhp�Y��`��sb+����IK�h�=�6{Ǚ:_���������ߍ����B�"@sMGK:�`P�Q��Ls��A,p|��{'�ڤW�/D?EWp�c��؊�o9M��
��M�'�c�{y�z��e�#�F�l<�B��]O��%۰O%��<r�e5C�f_��!>�ν���g��_��/gL��f�#�EgN()-#\$�\�Y���DB>'d�f��d?���@4�7h�
ǉ9���x�5�������:V19q���WxQ $���%��56��	�2��ea$�E����Ғ	�tlRh��`	d-f�Ԓu���:&�h�S�3��я.˨��v�ٜ���j$cT��	�$7~U4��Βy���&��=���Y��!1b({�o��rz3Pǌ�:֦�<G4�R<E�e�̼螪oJ�e�=��{�ތG���#��Mx}I�����G���1[g���X��p��ѥ,ߋu�e�&N��<.Y�WNH�k�|c?��M�
�t>�,�s|�2#b��-j)�������o?�ǘ�}�U�ˉ�V.f^��q�`x�9��K�!m'�������7�-�QMs�E�`λ�_Nz3
?�;�e�͊��~�]T$r�Ɗ/U��
}B^���c�k���~���7�jF�.l�g��^pr�3��+q#��)������{�{�H��C���c�L鈈�B��\�c���ġ��q���jh���@d^�Ѯii{���;p��e}w9��l�����YT�'_!ߚ;���¥HfH�+�2k�5�ASF�j�ʙ·P:{���s��	��d	��pT��!i����x~p󂭡�RS�R\o�"V�XLq/	@�U`,0�������""����*܍u�P�xC�|A7K�e#,�b�m��:��*�8�NB�������X��[���J汁w?���h��09qװ��~�g�(�5�׭�F�J���_�J���b��5Ƹr����z:P^��kϹI��\��7��������%��|�SB�/�[Q��"��ƚrK��T��(�R��T#����-K3uwUi�4_I®g����x��t�S$/�������v�"'V��c���)ʮl�R�Fp�I�xrQ'f$��[������X�%Z)	��t7^�RƄ��g��:_�ޘ�K��������.���*�|�!���K��s�?��Rl9g����fr��F���f��J�CrVZ��_�S���!�Q�̛��D'~�A����W�E�pP!.QC~:�/�y��$�c��3��4��֋��ULM��W0Q�v#�C/�B�9��q�=�݄	 S���E���}�AX��a��*� WMa��ə�qOu���EDO��k�ء��NF"|V1r�>�R�ʨ+1�T��@	'��x-x��ˏ�g�ea�{&z��6=O5���p1c���X+���cQ9bǆ�����dj���[���d-*b|Hvցޫ��i�zeG	{i�*.�P�a*`��!���]}߷NM:V�hR��~�
�v$|�RP����(����'�c{!��8�[z��!p`�����B��۟�֚�-T7!��0 ���A�Ԑ��@�$�9	��#��AV��ZO�TL�����N���V��@�2�x�M`�w����@T�'��B|�T��)��J��o��))��9)ӢD��s�a�!8t��le�%?'B��p���?�F씿��������_6_=UbkN��Mj��Y�d�_|�{1D99k6��Z8AM��ƪ�����rF�Aq�� MWZ��m'FM����;-��<|��t�mN��a��O߰�O����O�',���;_�h��u���sm��$W�S�HĊ��ԅsv�wث
�� ��2E��4���a��y��ܖ���䒺���x���X�>/�X������w;Q��kG��J�ի�q �6ǰ=��I�u��F$���س]8���3�F�j��)�/!ݲr��Ք��4��l��hgf����c�&�IK��6�!�Q0���x=��]=���,��d� ������0;����=��i�@w����sk).�sOvA�y��W��oh��6#��Mbۍ	Fm�����F�F�2��PK   �rZ,�_xU  �C     jsons/user_defined.json�[[o�F�+�-�Ý��o��t�ul�N�(E1ׄ�2�PR���ߏ��&)R�����Ky���;�e.�N�o�t����S^�0ݛ��y^��pF��|��[�����z���^��Ta�����9���"~(��p��M�җŢ*g�XM�k���x������4��Sʂ3���Hq���!�\QBqN��8�s_�7�U#��/r��Ac�� �AZ���2zN��*�)>�s铫����jY���M^�����:-��G��ff?��y�V�	�e}���m��Ճ�QZ��%��8	W�*:���r�����
a�\���
��������Z��̬��]���]M��%mX�{7���'�ǯ{aiV������emX9
�e�}/*o��Q��S�1�(����_�l���U-P�G���k}��JG��^L���Q�SL�o�mY�q�@�Aۢ�������%E����m��3���֓1x��AЫ��~�EᑰG���"�`69@Җ��p7����E�8�#�����"|,l�hG�ca�EK;����_hG�R#aM?jG��#Qu?j[c�����Q��d$��GmK�	cP���[l$j�C����D��]b$j��XG�#Q���:���
���Ic߮j�ۼ�d�7x
R�U��%�\3��q�rL;��]���X�K�o��&V���t��7櫆B��!�o��찳eSQ@+�����K�?����ay}��u-�>��n�\��e��&�������d�bYAa�zU� 5���G�"�����Q���i	uҪx����O����y�����U~}��E� �������ˬ��f��X\y�g�#�B>�(	�=q!Hk�W>�$k�L ȭ��`���Z)�S�ݿ�u�eUDY&k# �����,~ؐv��{xFz��6#ޢN��xB =�����f�m�o՛P�Aw��[x���Xj�|����d@�p��
j��*�$�˟/�pm�riK�/'o�y`.OQ"ceD!J�O�ٝ=���N���'oo�	���7��o7X~���Td$2䅰��X�g"RI��&I�'�<_.6h򑞂�:h�A��"5E.J��H!Y��g�	^i��xd��fZ�6�6�X��{�$�gHz��e����D4f}Sk���Mc��D�T�B�t	�����WJ�c�?O�\ He��^U����	ck��@��"�E�)���B	G��1Y�~/�B���iP���	E�����$%5	^�f���J5�R@`HS�!�	�i�(���O>z�vJ��*UI�WR���a�"*�T!#�A�� �Z��{)��l�!�5�%��Xi��
"*ᵦ��ϛi�g�U����|����D.y����)ͱ;݉�O)�#��_I�*fl륪hj�r��H�[�a����3�'���U���\.&��Uh��ar�W~��e���U���E��N:Ȏ�A[��I.�`cLI�r���u�ɑ���3���*���F��D��O4��$�9�1��4i���CFk��R�i���)e蝱o��y]�iN�8�L��f�pRL��wMC@��@�ta��l�n1���b�kkO���A����?G؞z�+�]��6�Ӱbŀ�V�s��)Y�0H��b�K�X���f�4R�ܿ�ڱ��@D��+x9���a��kA��j��� ���?�_���wy�j2����6+���c��r��[ӌ)�ɞ��&�j�����I=u���%�5�dZ��89�~��-}��z4�ǧ��� j{ ݌�?�ia��s~yp���ȵ�Z���D��Gw,�s�r���v&p��t�Ţ,��w�'�q~Cط	�9Ɉ��q"�N
���,�d96�[LU��=UgB�+��J�562-�	{�t� ���9�R�a��/c��2�A!�\|�E�^���<U��������tА�7y��ұ�}�w$#L|d�p��Jrqu*0����WD�p���'��r��t� �9C5b>F�sA
|dX2�N�`��;���;���;���;���;���;��{�<�RN^-���7�g����p1Q�G���0\�zg�C6Pm�^
3�[Dd�����$��*� a4S_�
!2"U���KDf�t{_B0�S����?�ٓ���-@p�Z�$+x14W�ӱS]k�S�Z&G��s	n�^G���pU�[]ۮN�����������P��e8!X{���~br�rp&�>���Q�y�D��`�47H�DQ�[O�掷��RSh��0:�r�4�c�Q���#�͔�W���ֿm�$'�h\87<3|0�m<��	�i�i6#�n��T�L�a����5!nM 6�I5��>�3Flm�܂(�I����y,��S��)c���r��UJ"Ǭ��@��(�)�|�(F�	V#gA<J��vy̴��媽��e�*�������,1AC0�9�^@(,3��N���m=���tr�՞��[u��r�(�l�m�j��V��洩ܚ�Q��L��W?�\��joꕷ7�e���D��P�"bN1�4.���X���̖K�C]sDi�Ղ:�YC���_m�S��� +x�����Ӓ�=� �4�W�@n��A6��)��Xy���p�[{ё�5�m=��������mN@�m).�G���fC&=�#�B<(����V�n�&�,����g^&��1�Ƅ _��E�
�XD�Jd�!uÆ��<dM�GH,I�gRΜ�_CF3<P��u	Mg�h�����zjĞʔ�ٖ'e(��)��2�Yb�s2�n��B������J���<<�"����9����z�|���a�,#�JH&��]����PK
   �rZrr���=  ��                  cirkitFile.jsonPK
   �}rZ�$&VAS }d /             �=  images/6227b039-7cc5-4ac4-8a39-c32f35a7f912.pngPK
   r}rZר� �* /             �� images/731a9da8-b9b1-4e67-98b9-c038a7318a47.pngPK
   G�rZ�SIM7#  2#  /             � images/7346828c-be13-4248-836b-104e84d3cd43.pngPK
   ��rZ�c^��  �  /             p� images/7daa3674-301d-466b-aa13-7b9309bd01d6.pngPK
   �rZ��p� �� /             � images/7e81f6ad-0912-4ff6-bfc6-e58bb7840941.pngPK
   G�rZ�mg��S �S /             Ҵ images/84f81591-1534-4849-82f2-ec60ac1f84b4.pngPK
   �rZ�1.:�  )  /             		 images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.pngPK
   �rZ?S��� 2� /             "(	 images/99226213-8268-43da-ade8-d9d07cfcec9f.pngPK
   �}rZ"1^F�� Ho /               images/a027fa6b-1779-4bc7-b1bd-261c8096f986.pngPK
   �}rZ����  �  /             � images/a36c4c40-5e17-4d78-b145-5ddca5d02051.pngPK
   �}rZ������  ��  /             B� images/a4634dc7-be5e-40a8-852b-d0b700abe16e.pngPK
   �rZ$�8�l  �  /             G� images/aa130aff-16e6-4627-9689-819d55b5861f.pngPK
   �rZ���7z  �  /              � images/be8de2bb-09ef-440a-a2d8-19619bf9d0dd.pngPK
   �rZ6e�b�  �  /             �� images/c0cd0a79-4e96-4647-8bb3-400a2b193618.pngPK
   �rZ;mLF   P   /             �� images/c560fc9b-7045-4fe6-9a6e-de67d6663603.pngPK
   �rZ$7h�!  �!  /             8 images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   �}rZ��@�/  �/  /             {0 images/c6f01788-a49f-442a-a7cf-1585482f8cc6.pngPK
   r}rZ���O!	 � /             \` images/cbf232a7-7072-4b1f-a35a-352dd9a3bcf3.pngPK
   �rZ�^X�� j( /             �i images/cfd750a9-6fd4-4ac0-902f-08baa65eb73b.pngPK
   �rZ�GDU7� �� /             � images/d628d844-ce42-4e82-be63-f5fdfa438334.pngPK
   ��rZ A��?5 �J /             ol images/e0d6f4e0-adc9-461d-95f3-67e9d6b55837.pngPK
   �rZP��/�  ǽ  /             �� images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   �rZF���?� Q� /             MT images/f590943e-678c-44eb-a174-3243ba5f3820.pngPK
   �}rZ��g  n  /             �� images/f636b928-3cee-4f31-b55b-93d56e3d5b88.pngPK
   �rZ,�_xU  �C               �� jsons/user_defined.jsonPK      :	  
    